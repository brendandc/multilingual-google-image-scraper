ab	ab
abba	abba
abbas	abbas
abbey	abbey
abc	abc	abc (swedish news program)
abort	abortion
aborter	abortions
about	about
abraham	abraham
absint	absinthe
absolut	absolute; total	absolute
absoluta	absolute
absolution	absolution
absorberas	(gets) absorbed
abstrakta	abstract
abu	abu
ac	ac
academy	academy
acceptera	accept
accepterad	acceptable
accepterade	accepted
accepterar	accepts	accept
accepterat	accepted
acdc	ac/dc
action	action
ad	ad
adam	adam
adams	adams
adeln	nobility
adhd	adhd
adjektiv	adjective	adjectives
administration	administration
administrationen	administration
administrativ	administration	administrative
administrativa	administrative	administative
administrativt	administrative	administratively
adolf	adolf
adolfs	adolf's
adrian	adrian
advokat	lawyer
af	of (old swedish)
affärer	business
afghanistan	afghanistan
africa	africa
afrika	africa
afrikaner	africans
afrikansk	african
afrikanska	african
afrikas	africa's	africas
afrodite	afrodite
aftonbladet	aftonbladet	the evening paper
age	age
agent	agent
agera	act
agerande	acting	behavior
aggressiv	aggressive
agnes	agnes
agnetha	agnetha
agnosticism	agnosticism
agnostiker	agnostic	agnostics
ahmed	ahmed
aids	aids
aik	aik
airlines	airlines
airport	airport
ajax	ajax
akademi	academy
akademien	the academy	academy
akademiens	the academy's
akademisk	academical	academic
akademiska	academical	academic
akc	akc
akon	akon
akondroplasi	achondroplasia
aktiebolag	companies	limited company; joint-stock company	stock company
aktier	stock
aktiv	active
aktiva	active
aktivitet	activity
aktiviteten	activity
aktiviteter	activities
aktivt	actively
aktuell	current
aktuella	current
aktuellt	current	relevant
aktörer	players	actors
akut	acute	urgent
al	alder
alan	alan
alaska	alaska
albaner	albanians
albanien	albania
albanska	albanian
albert	albert
album	album
albumen	the albums	albums
albumet	album
albumets	album's
alces	alces
aldrig	never
ale	ale
alex	alex
alexander	alexander
alexanders	alexanders	alexander's
alexandra	alexandra
alexandria	alexandria
alf	alf
alfa	alpha
alfabet	alphabets	alphabet
alfabetet	alphabet	the alphabet
alfabetisk	alphabetical
alfred	alfred
alger	algaes
algeriet	algeria
ali	ali
alice	alice
alkohol	alcohol
alkoholer	alcohols
alla	all	everyone
allan	allan
alldeles	completely	altogether
allen	allen
allians	alliance
alliansen	the alliance
allierad	allied	ally
allierade	allied
allierades	allied's	allied
allmän	general
allmänhet	in general	general
allmänheten	public	general public
allmänna	general
allmänt	commonly	generally; public
allra	very	most	-most; most
alls	all
allsvenskan	allsvenskan
allt	all
alltför	all too	exessive
alltid	always
allting	everything
alltjämt	remains
alltmer	increasingly	more and more
alltsedan	even since	since
alltså	so	therefore	really
allvar	earnest
allvarlig	serious
allvarliga	serious
allvarligt	serious
alperna	alps	the alps
alqaida	al-qaida	al-qaeda
alternativ	alternative
alternativa	alternative
alternativt	alternatively	alternative
aluminium	aluminum
am	am
amazonas	the amazon rainforest	amazonas
ambassad	embassy
ambitioner	ambitions
america	america
american	american
amerika	america
amerikanen	american	the american
amerikaner	american	americans
amerikanerna	the americans
amerikansk	american
amerikanska	american	u.s.
amerikanske	american	the american
amerikanskt	american
amerikas	america
amfetamin	amphetamine
aminosyra	amino acid
aminosyror	amino acids
ammoniak	ammonia
amsterdam	amsterdam
amy	amy
ana	feel
analsex	anal sex
analys	analysis
analytisk	analytical
analytiska	analytical
anarkism	anarchism
anarkismen	the anarkism	anarchism
anarkister	anarchists
anarkistiska	anarchistic	anarchist
anatolien	anatolia
anatomi	anatomy
anc	anc
anda	spirit
andas	breath
ande	of	spirit
andel	share
andelen	share	the share	the proportion
anden	the holy spirit
anderna	andes	the andes
anders	anders
andersson	andersson
anderssons	anderssons	andersson's
andlig	spiritual	spirtual
andliga	spiritual
andra	second	other
andras	others
andre	other
andreas	andreas
andres	andres	other's
andrew	andrew
andré	andre
andy	andy
anfall	attack
anfalla	attack
anfallet	the attack	attack
anfield	anfield
anföll	attacked
ange	set	name
angeles	angeles
angelina	angelina
angels	angels
anger	indicates	gives
anges	mention	is put at	specified
anglosaxiska	anglo-saxon
angola	angola
angrepp	attack
angränsande	adjoining
angående	concerning	reference
anhängare	followers	supporters
anhöriga	relatives	kin
animerade	animated
anka	anka	duck
anklagade	accused
anklagades	accused
anklagats	accused
anklagelser	allegations	accusations
anknytning	tie	link
ankomst	arrival
anlades	were built
anledning	reason
anledningar	reasons
anledningarna	reasons	the reasons
anledningen	reason
anläggningar	facilities
anlände	arrived
anländer	arrive	arrives
anna	anna
annan	another
annars	else
annat	other	other; another
anne	anne
annekterade	annexed
annika	annika
annorlunda	different
anor	ancestry	lineage; ancestry
anordnas	provided	arranged
anorektiker	anorectics	anorectic
anorexia	anorexia
another	another
anpassa	adjust	adapt
anpassade	custom
anpassat	adapted
anpassning	adaption
anser	view	believes
anses	deemed; regarded
ansetts	regarded	regarded; viewed (as)
ansikte	face
ansiktet	face
ansluta	join	connect
ansluter	connects
anslutna	affiliated
anslutning	connection
anslöt	joined
anspråk	claim	claims
ansträngningar	effort
anställd	employed	hired
anställda	employed
ansvar	responsibilities	responsibility
ansvarar	charge
ansvaret	responsibility	the responsiblity
ansvarig	charge
ansvariga	charge
ansåg	thought	considered	found
ansågs	was	seemed
ansökte	applied
anta	assume	adopting	assume; adopt
antagit	presumed
antagits	adoption	adopted
antagligen	ligands presumably	probably	presumably
antal	number of	number
antalet	number	the number
antar	adopting	suppose
antarktis	antarctica
antarktiska	antarctic
antas	is required	expected (to)
anteckningar	notes
anthony	anthony
antika	ancient
antiken	the ancient world
antikens	the ancient's	ancient
antingen	presumably	either
antisemitiska	antisemetic	antisemitic	anti-semitic
antisemitism	antisemitism
antisemitismen	antisemitism	anti-semitism
antog	adopted
antogs	was assumed
antoinette	antoinette
antonio	antonio
antropogen	anthropogeny	an anthropogenic	antropog	antropogenic	man-made	anthropogenic
antyder	indicates
anus	ass	anus
använda	using
användande	use	use; usage
användandet	usage	use
användare	users
användaren	the user	user
användas	used
användbar	useful
användbara	usable	useful
använder	using	uses
användes	was used	used
användning	use	use; usage
användningen	use	the use
användningsområden	possible use	applications
används	use	used
använt	used
använts	was used	used
apartheid	apartheid
apollo	apollo
april	april
ar	is
arab	arab
arabemiraten	united arab emirates	uae	the arab emirate
araber	arabs
araberna	arabs
arabisk	arabic
arabiska	arabic	arabian
arabvärlden	the arab world	arab world
arbeta	work	working
arbetade	worked
arbetar	work	works
arbetare	workers
arbetarklassen	working class	the working class
arbetat	worked
arbete	work	work; labor
arbeten	works
arbetet	work	the work
arbetsgivare	employers
arbetsgivaren	employer
arbetskraft	workforce	labor
arbetslöshet	unemployment	unemplyment
arbetslösheten	unemployment
arbetsplats	workplace
area	area
arean	the area	the space
arena	arena
arenan	arena	the arena
arg	angry
argentina	argentina
argument	argument	arguments
aristokratin	the aristocraty	aristocracy
aristoteles	aristoteles	aristotle
arkeologiska	archaeological
arkitekt	architect
arkitekten	the architect
arkitekter	architects
arkitektur	architecture
arkitekturen	the architecture	architecture
arkiv	archive	archives
arlanda	arlanda
arm	arm
armar	arms
armenien	armenian
armeniska	armenian
army	army
armé	army
arméer	army
arméerna	armies
armén	the army
arméns	the army's	army's
arnold	arnold
arrangemang	arrangement
arrangeras	(is) arranged	arrange
arresterades	was arrested
arsenal	arsenal
art	kind	art
arten	species
arter	species
arterna	the species	species
arternas	the species
arthur	arthur
artikel	article
artikeln	the article
artiklar	items
artist	artist
artisten	the artist
artister	performers	artists
artisterna	aristerna
arton	18	eighteen
arvet	the inheritance
arvid	arvid
asiatiska	asiatic	asian
asien	asia
aspekt	aspect
aspekter	aspects
aspergers	downs syndrome	aspergers
assistent	assistant
assisterande	assistant	assisted
assyriska	assyrian
asterix	asterix
asteroidbältet	the asteroid belt
asteroider	astroids	asteroids
aston	överraska, undra	aston
astrid	astrid
astronomer	astronomers	astronomer
astronomi	astronomy
astronomin	the astronomy
astronomiska	astronomical
ateism	atheism
ateist	atheist
ateister	atheists
aten	athens
atlanta	atlanta
atlanten	atlantic	the atlantic ocean
atlas	atlas
atmosfär	atmosphere
atmosfären	the atmosphere
atom	atomic	atom
atombomben	the nuclear bomb
atombomberna	atom bombs	the nuclear bombs	atomic bomb
atomer	atoms
atomkärnor	nuclei	nuclear particles	atomic cores
att	to	that
attacken	the attack
attacker	attacks	assaults
attackerna	attacks	the attacks	attack
august	august
augusti	august
auktoritet	authority
auktoritära	authoritarian
auschwitz	auschwitz
austin	austin
australia	australia
australian	australian
australien	australian	australia
australiens	australia's
australiska	australian
autism	autism
automatiskt	automatic
autonom	independent	autonomic
autonoma	autonomous	autonomic
autonomi	autonomy
av	of
avalanche	avalanche
avancerad	advanced
avancerade	advanced
avbrott	break
avbryta	cancel
avbröts	canceled	interrupted
avel	breeding	breed
avfall	waste
avgick	resigned	retired
avgå	resign
avgör	decides
avgöra	determine	decide
avgörande	settling	decisive
avgörs	determined	decided	is determined
avhandling	treatise	thesis
avkomma	progeny	offspring
avled	deceased	died
avlidit	perished
avlidna	diseased	deceased	the perished
avlägsna	remove
avrättades	was executed	executed
avrättning	execution
avrättningar	execution	executions
avrättningen	execution	the execution
avsaknad	absence
avsaknaden	absence
avsattes	deposited	dismissed
avsedd	intended
avsedda	intended	aimed
avseende	regard
avseenden	regard
avser	regards	regard
avses	regard	referred
avsett	regard	intended
avsevärt	substantially	considerably
avsikt	intention
avsikten	intention	purpose
avskaffa	abolish
avskaffade	abolished
avskaffades	was abolished	abolished
avskaffande	abolition	abolishment
avskaffandet	abolition	abolishment
avsluta	finish	exit
avslutade	ended	finished
avslutades	ended; concluded
avslutas	close	ends
avslutat	completed	finished
avslöjade	revealed
avsnitt	part	episode
avsnitten	the episodes	chapters
avsnittet	episode
avstå	desist	refrain
avstånd	distance
avståndet	the distance
avsätta	unseat
avsåg	meant	mean
avtal	agreement; deal	contract
avtalet	the treaty	the contract	agreement
avtar	declines
avvikande	different	deviant; divergent; different
avvikelser	deviations	derivations
avvisade	rejected
avvisar	reject
awards	awards
axel	axel
axelmakterna	the axis	axis
axl	axl
azerbajdzjan	azerbaijan
azidgrupp	azido group	azid group	azide group	azide	amide
b	b
babylon	babylonia	babylon
bad	bath
bagge	ram
bahamas	bahamas
baháulláh	bahullah
baháí	bahá'í
baker	baker
bakgrund	background
bakom	behind
bakterier	bacteria
bakåt	backwards	reverse
balans	balance
balansen	balance	the balance
balkan	the balkans
balkanhalvön	balkan peninsula
baltikum	the baltics	baltics
baltimore	baltimore
baltiska	baltic
bana	course
banan	the track	banana
banbrytande	groundbreaking
band	band	tape
banden	bander	the bound
bandet	band
bandets	the bands	band
bandmedlemmar	band members
bandmedlemmarna	band members
bank	bank
banker	banks
banor	paths	line
baptism	baptist	bapist faith	baptist faith	baptists	baptism	döpare
bar	bar
bara	only
barack	barracks
barbro	barbro
barcelona	barcelona
barcelonas	barcelona's
barndom	childhood
barnen	children
barnens	childrens
barnet	child
barnets	the childs	the child's
barney	barney
barns	childrens	children	child
baron	baron
barrett	barett	barrett
barry	barry
bars	carried
bart	offense	bart
bas	base
basen	became	the base	base
baser	bases
baserad	based
baserade	based
baserar	base	based
baseras	based	bases	based on
baserat	based
basis	basis
basist	bassist
basisten	basist	the basist
basket	basketball
batman	batman
bay	bay
bayern	bayern
bbc	bbc
be	be
beatles	beatles
bebott	inhabit	inhabited
bebyggelse	settlement	settlements	habitation
bebyggelsen	settlement
beck	beck
beckham	beckham
bedrev	conducted	managed
bedriva	carry	prosecute
bedriver	manage	operate
bedrivs	conducted
bedöma	judge; decide
bedöms	judged	evaluated
beethoven	beethoven
befann	located	found
befinna	be
befinner	is	placed; situated; positioned; are
befintliga	existing
befogenhet	warrant	authority	authorization
befogenheter	authorities	powers
befolkade	inhabitated	populated
befolkning	population
befolkningen	the population
befolkningens	population's
befolkningstillväxt	befolkningstillvaxt	population growth
befolkningstillväxten	population growth	the population growth	the growth of population
befolkningstäthet	population density
befolkningstätheten	population density	state of the population
befolkningsutveckling	population development	population growth
befruktning	conception	fertilization	conceptions	fertilizing	fertilisation	insemination	impregnation	monograph
befäl	command
befälet	the command
befälhavare	commander
begav	went	traveled	went (to)
begick	commited	committed
begravd	buried
begravdes	buried
begravning	funeral
begrepp	term	concept
begreppen	the concepts	the terms
begreppet	term	concept
begränsa	limit
begränsad	limited	restricted
begränsade	restricted	limiting
begränsar	limit	limits
begränsas	limited	(gets) limited	begransas
begränsat	restricted	limited
begränsningar	limitations
begär	requests
begäran	request
begärde	called	demanded
begå	commit
begår	commit	commits
begått	committed	comitted
behandla	treatment
behandlade	was treated	treated
behandlades	treated
behandlar	treats	treat
behandlas	treated
behandling	treatment
behandlingar	treatments
behandlingen	the treatment	the treament	treatment
behov	necessary
behovet	need	the need
behålla	keep
behåller	retain	keeps
behöll	kept
behöva	need
behövde	needed
behövdes	required
behöver	need
behövs	required	is needed
bekant	known	acquaintance
bekostnad	expense
bekräftade	confirmed
bekräftades	confirmed	was confirmed
bekräftar	confirms
bekräftat	confirmed
bekämpa	prevent	combat; fight	fight
belagt	coated
belgien	belgium
belgiens	belgium's
belgiska	belgian
belgrad	belgrade
bell	bell
bella	bella
belopp	amounts	amount	sum
belägen	located	situated
beläget	located	base
belägg	evidence
belägna	located
belönades	rewarded	awarded
bemärkelse	meaning	sense
ben	bone
benen	legs
benfica	benfica
bengt	bengt
bengtsson	bengtsson
benny	benny
bensin	gasoline
benämnas	named	entitle	entitled
benämning	term	name
benämningar	terms	names
benämningen	the designation	the name	label
benämns	designated	is mentioned
beordrade	commanded	ordered
ber	asks
beredd	ready (to)	prepared
berg	mountain(-s)	mountain
bergarter	rock types	minerals	rocks
bergen	mountain
berger	berger
berget	mount	the mountain
bergman	bergman
bergmans	bergman's	bergmans
bergqvist	bergqvist
bergskedjan	mountain range	the mountain group
bergskedjor	mountain ranges
berlin	berlin
berlinmuren	berlin wall	the berlin wall
berlins	berlin	berlin's
bernadotte	bernadotte
bernhard	bernhard
bero	depend
berodde	was	depended
beroende	dependent	depending
beroendeframkallande	addictive
beror	is
bertil	bertil
beräkna	calculate
beräknades	estimated
beräknar	computes	values
beräknas	estimated
beräkningar	calculations
berätta	tell
berättade	told
berättar	tells
berättas	(as) told	is told	told
berättat	told
berättelse	tale	story
berättelsen	story	the story
berättelser	tales	stories
berättelserna	the stories	tales; stories
berömd	famous
berömda	famous
berömt	famous	praised
berör	affect	concerns
besegra	defeat
besegrade	defeated
besegrades	defeated
besegrat	defeated
besittning	dominion	possess
besittningar	holdings
beskrev	depicted	described
beskrevs	was described	described
beskriva	describe
beskrivas	described	be described
beskriver	describes
beskrivit	described
beskrivits	described
beskrivning	description
beskrivningar	description	descriptions
beskrivningen	description
beskrivs	described
beskydd	protection
beskyddare	protector	patron
beslut	decision
beslutade	decided
beslutar	decides
beslutat	decided
besluten	decisions
beslutet	the decision
besläktade	related
besläktat	related to	related
beslöt	decided
besserwisser	pundit	smartass	bewiseacre	exact: better knower; equivalent: know-it-all	know-all	know-it-all	know it all	besserwisser	wiseacre
best	best
bestod	was
bestämd	fixed
bestämde	determined	chose
bestämdes	was decided	decided	was determined
bestämma	determining	decide
bestämmelser	regulations	measures
bestämmer	decide
bestäms	is decided
bestämt	decided
bestå	consists	exist	comprise
bestående	comprising	lasting
beståndsdelar	constituents	elements
består	consists of	exists
besättningen	crew
besök	visit
besöka	visit
besökare	visitors
besöker	visits
besökt	visited
besökte	visited
bet	bit
beta	beta	graze
betala	pay
betalade	payed	paid
betalar	pay
betalt	charge
beteckna	denote
betecknar	represent	denotes
betecknas	denote	labelled	designate
beteckning	label
beteckningen	the label	designation.........	designation
beteende	behaviour	behavior
beteenden	behavior
betonade	emphasized
betonar	stress	emphasize
betoning	stress
betrakta	view; regard
betraktade	considered
betraktades	considered	regarded
betraktar	regard
betraktas	considered
betraktats	considered	(been) viewed
betyda	mean
betydande	important
betydde	meant	ment
betydelse	significance
betydelsefull	meningful	significant
betydelsefulla	significant
betydelsen	the meaning	significance
betydelser	meanings
betyder	means
betydligt	considerably	significant
betyg	grades
bevara	preserve
bevarad	kept	preserved
bevarade	preserved
bevaras	are protected
bevarat	preserve	preserved
bevarats	protected	preserved
bevis	certificate	evidence
bevisa	prove
beväpnade	armed
beyoncé	beyonce	beyoncé
bibel	bible	bilble
bibeln	bible
bibelns	the bibel's	the bible's	bible
bibliografi	bibliography
bibliotek	library
bibliska	biblican
bidra	contribute
bidrag	contribution
bidragande	contributors
bidragen	the contributions	contributions
bidraget	grant
bidragit	contributed
bidrar	contributes
bidrog	contributed
big	big
bil	car
bilar	cars
bilbo	bilbo
bild	picture
bilda	form
bildade	formed
bildades	founded	was formed
bildande	founding	formation
bildandet	establishment
bildar	serves as	form
bildas	formed; made up (of)	formed
bildat	formed
bildats	had formed	created
bilden	the image
bilder	pictures
bilderna	the pictures
bildning	education	form	learning
bildt	bildt
bilen	the car	car
billboardlistan	bilboardlist
billiga	cheap
billy	billy
bilmärke	car make	make of car
binda	bind	tying
bindande	binding
binder	tie	bind
binds	bound	(is) bound
bioetik	bio ethics	bioethic	bioethics
biogeografi	biogeography	biogegraphy
biografen	the cinema	movie theater
biografer	movie theaters	movie theaters; cinemas	cinemas
biografi	biography
biologi	biology
biologisk	biological
biologiska	biological
bipolär	bipolar
bipolära	bipolar
birger	birger
birgitta	birgitta
birk	birk
birmingham	birmingham
biskop	bishop
biskopen	bishop	the bishop
bistånd	aid
bit	piece
bitar	pieces
biträdande	assistant	assisting
bitter	bitter
bjöd	invited	offered
björn	björn
bl	short of "bland" - in the context: bl. a (bland annat) = among others
bla	blah	among others
black	black
blad	leaves	leaf
blanc	blanc
bland	inter	including
blanda	mix
blandad	mixed
blandade	mixed
blandas	mixed	mixes
blandat	mixed
blandning	mix	mixture
blekinge	blekinge
blev	became
bli	become
blind	blind	bank
blir	become
blivande	prospective	future	to be
blivit	become
block	block
blod	blood
blodet	the blood	blood
blodiga	bloody
blodkroppar	corpuscle
blodtryck	blood pressure
blodtrycket	the blood pressure	blood pressure
blogg	blog
bloggar	blogs
blommor	flowers
blomstrade	flourished
blott	merely	mere
blue	blue
blues	blues
bly	led	lead
bläckpenna	pen	ball point pen	ink pen	ball point pen; pen	black pen	quill
blå	blue	blah
blåser	blowing
blått	blue
blåvitt	blåvitt	bluewhite	blue and white
bmi	bmi
bnp	gdp	gnp
bob	bob
bobby	bobby
bodde	lived
boende	resident
bojkott	boycott
bok	book
boken	paper	the book
bokförlaget	bokförlaget	publisher	publishing house
bokstav	letter
bokstaven	the letter	character
bokstäver	letters
bokstäverna	the letters
bolag	company
bolaget	the company
bolagets	company's	the corporation's
bolivia	bolivia
bolivianska	bolivian
bolivias	bolivia's
bollen	the ball	ball
bolsjevikerna	the bolsheviks
bolt	bolt
bomb	bomb
bomben	the bomb
bomber	bombs
bomull	cotton
bon	bon
bonaparte	bonaparte
bond	bond
bonde	farmer
bonniers	bonnier's	bonniers
book	book
bor	lives
bord	table
borde	should
bordet	the table
borg	castle	tower
borgen	castle	bail	the castle
borgerliga	conservative
borgmästare	mayor
boris	boris
born	born
borrelia	borrelia	borreliosis
bort	away	remove
borta	gone	away
bortgång	passing
bortom	beyond
bortsett	except
bosatt	resident	lived
bosatta	residents	settled
bosatte	settled
bosnien	bosnia
bosnienhercegovina	bosnia-hercegovina
bostad	lodge
bostadsområden	residential	housing	residential areas
boston	boston
bostäder	residences	housing
bosättare	settlers
bosättningar	settlements	bosattningar
bott	lived in
botten	the base	bottom
bowie	bowie
boxning	boxing	boxing; pugilism
boy	boy
bra	good
brad	brad
brand	fire
branden	the fire
brandenburg	brandenburg
brasilianska	brasilian
brasilien	brazil
brasiliens	brazil's
breaking	breaking
bred	broad
breda	broad	qual o curso que você está estudando	wide
bredare	wider
breddgraden	latitude	parallel
bredvid	beside	next to
brev	letter
brevet	the letter
brian	brian
bridge	bridge
brinnande	burning
brinner	on fire
brist	non	failure; lack of
bristande	wanting	lack
bristen	lack of
brister	inabilities
brita	brita
britannica	britannica
british	british
britney	britney
britter	britons
britterna	british	the brits
brittisk	british
brittiska	british
brittiske	british
brittiskt	brittish	british
bro	bridge
broar	bridges
broder	brother
brodern	the brother
bron	the bridge
brons	bronze
bronsåldern	bronze age	the bronze age
bronx	bronx	the bronx
brooke	brooke
brooklyn	brooklyn
bror	brother
brother	brother
brott	breach	crimes	crime
brottet	offense	the crime	the crime; offense; infraction; transgression
brottslighet	criminality	crime
brottslingar	criminals
brown	brown
bruce	bruce
bruk	use
brukade	used to	used
brukar	usually	used to
bruket	the use
brushane	ruff
brutit	cut; break	broken
bruttonationalprodukt	bnp
bryssel	brussels
bryta	break
bryter	breaks	breaking; violating
bryts	breaks
bränder	fires
brändes	burned	burnt
brännvin	schnaps	aquavit
bränsle	fuel
bränslen	fuel
bråk	brawl; fight	fights
bröd	bread
bröder	brothers
bröderna	brothers	the brothers
bröllop	brollop	wedding
bröllopet	the wedding
bröstet	chest; breast	breast
bröt	brot	broke
bröts	was fractured	broke
bud	bid	message
budapest	budapest
buddha	buddha
buddhas	buddha's	buddhas
buddhism	buddhism
buddhismen	buddism
buddhister	budhists	buddhists
buddhistiska	buddhistic	buddhist
buddy	buddy
budet	the bid	the commandment
budget	budget
budgeten	budget	the budget
budskap	message
budskapet	message	the  message
bulgarien	bulgaria
bulgariens	bulgaria	bulgaria's
bulgariska	bulgarian
bundna	bound	tied
bunny	bunny
burj	burj
burma	burma
burr	burr
burton	burton
burundi	burundi
bush	bush
bushadministrationen	the bushadministration	the bush administration	bush administration
bushs	bush's
buss	bus
bussar	bus
butiker	shops
by	village
byar	villages
bygga	build
byggandet	the building
byggas	build
byggd	built
byggda	constructed
byggde	built	built, founded (on)
byggdes	was built
bygger	based	(is) building (on)
bygget	the construction	construction
byggnad	building
byggnaden	building	the building
byggnader	buildings	structures
byggnaderna	buildings	the buildings
byggnadsverk	building	edifice
byggs	building	under construction
byggt	built
byggts	built
byn	village
byrå	its section	agency	bureau	office
bysantinska	byzantine
byta	switch	change	trade
byte	change of	bytes
byten	byte
byter	changes	exchanges
bytet	the exchange	change
byts	replaced
bytt	traded	switched
bytte	changed	swapped
byttes	changed	was exchanged
byxor	pants
bägge	both
bär	carryng	here	berries
bära	carry	mean
bärande	wearing	leading	fundamental; wearing; supportive
bäst	best
bästa	the best	best
bäste	best
bättre	better
båda	both
både	both
bål	prom	torso
båt	boat
båtar	boats
båten	the boat	boat
böcker	books
böckerna	books
böhmen	bohemia
bön	nests	prayer
bönder	farmers
bönderna	the farmers	farmers
bönor	beans
bönorna	beans
bör	live	should
bördiga	fertile
börja	start
började	started	began
början	beginning
börjar	starts
börjat	started	begun
börje	borje
ca	cirka	approximately
caesar	caesar
caesars	caesars
café	coffeehouse	café
california	california
calle	calle
cambridge	cambridge
camp	camp
campus	campus
can	can
canada	canada
canadian	canadian
canaria	canaria
cancer	cancer
cannabis	cannabis
cant	cant
capita	capita
capitol	capitol
carl	carl
carlo	carlo
carlos	carlos
carlsson	carlsson
carola	carola
carolina	carolina
carter	carter
cash	cash
casino	casino
castro	castro
cd	cd
cecilia	cecilia
cell	cell
cellen	cell	the cell
cellens	the cell's	cell's
celler	cells
cellerna	cells	the cells
census	census
center	center
centra	center
central	central
centrala	central
centralamerika	central america
centralasien	central asia
centralbanken	centralbank	central bank
centraleuropa	central europe
centralort	central city	regional centre
centralorter	regional centers	centers
centralstation	central station
centralt	central
centre	centre
centrum	center
champagne	champagne
chandler	chandler
channel	channel
chans	chance	chanse
chansen	chance
chaplin	chaplin
charles	charles
charlie	charlie
charlotte	charlotte
chefen	commendant; commander
chelsea	chelsea
chi	chi
chicago	chicago
chile	chile
chiles	chiles	chile's
chili	chili
choice	choice
choklad	chocolate
chokladen	the chocolate
chris	chris
christer	christer
christian	christian
christina	christina
chrusjtjov	chrusjtjov
church	church
churchill	churchill
cia	cia
cirka	about	approximately
cirkel	circular
citat	quote
city	city
civil	civil	civilian
civila	civil
civilbefolkningen	civilian population	the civilian population	civilians
civilisationen	civilization
civilisationer	civilizations
claes	claes
claude	claude
cliff	cliff
clinton	clinton
club	club
cobain	cobain
cocacola	coca cola	coca-cola
cohen	cohen - it's a name	cohen
coldplay	coldplay
colin	colin
colombia	colombia
colombo	colombo
colorado	colorado
colosseum	colosseum
columbia	columbia	colombia
columbus	columbus
come	come
comeback	comeback
comet	comet
cosa	cosa
costa	costa
counterstrike	counterstrike
country	country
county	county
cover	cover
craig	craig
crazy	crazy
crick	crick
cricket	cricket
criss	criss
cruz	cruz
crüe	crüe
cupen	the cup
cykel	bicycle
cykeln	there are two meanings in the context - cycle and bicycle	cycle
cyklar	bicycles	bikes
cypern	cyprus
cyrus	cyrus
da	da
dag	dag	day
dagar	says	days
dagarna	the days
dagars	day's	days
dagbladet	daily paper	dagbladet
dagbok	diary
dagen	day
dagens	current	todays
dagliga	daily
dagligen	daily
dagligt	daily
dags	time
dagsläget	present situation	current situation
dahlén	dahlén
dahléns	dahlens	dahlén's
dalar	valleys
dalarna	dalarna
dalí	dali
dam	dam	lady
damer	ladies
dancehall	dance hall
daniel	daniel
danmark	denmark
danmarks	denmark's
danny	danny
dans	dance
dansk	danish
danska	danish
danske	danish
dark	dark
darwin	darwin
darwins	darwins
das	das
data	data
dateras	dates
dator	computer
datorer	pc
datorn	the computer
datorspel	video game	computer game
datum	date
dave	dave
david	david
davis	davis
day	day
de	the	they
debatt	debate
debatten	the debate
debatter	debates
debut	debut
debutalbum	debut album
debutalbumet	the debut-album	debut album
debuterade	debut	debuted
december	december
decennier	decades
decennierna	decades	the decades
decenniet	decade
decennium	decade
deep	deep
define	define
definiera	define
definierade	defined
definierar	defines
definieras	is defined	defines
definierat	defined
definition	definition
definitionen	definition	the definition
definitioner	definitions
definitivt	unavoidable	definitely
deklarerade	declared
del	part
dela	divide	dividing
delad	shared	divided
delade	divided	split
delades	shared	divided	split
delar	proportions	parts
delarna	the parts	parts
delas	shared	divided
delat	divided
delats	divided	been awarded
delen	part
delhi	delhi
delning	division	pitch
delningen	division	pitch
dels	and	both	partly
delstat	state
delstaten	land	the state
delstater	states
delstaterna	states
delta	participate
deltagande	participation
deltagare	contestant	participiant
deltagarna	the participants	participants
deltagit	participated
deltar	participates
deltog	participated
delvis	partly	partial	partially
dem	those
demens	dementia
demo	demo
demografi	demographics	demography
demografiska	demographic	demographical
demokrati	democracy
demokratier	democracies
demokratin	the democracy	democracy
demokratisk	democratic
demokratiska	democratic
demokratiskt	democratic
demonstrationer	demonstrations
den	it
denna	that
denne	that he	he
dennes	his
dennis	dennis
densamma	the same	same
densitet	density
densiteten	density
departement	department
depolarisering	depolarisation	de-polarizing	depolarization
depp	depp
depression	depression
depressionen	the depression	depression
depressioner	recessions	depressions
der	where	german word
deras	their
derivata	derivative
derivatan	the derivative
derivator	derivative	derivatives
design	design
desmond	desmond
dess	then	its
dessa	these
dessförinnan	before (that)
dessutom	moreover	furthermore	furthermore; moreover, additionally; likewise
desto	ever
det	it	dent
detalj	detail
detaljer	details
detroit	detroit
detsamma	the same	same
detta	this
deuterium	deuterium
development	development
diabetes	diabetes
diagnos	diagnostics
diagnosen	diagnosis	the diagnose
diagnoser	diagnoses
dialekt	dialect
dialekter	dialects
dialekterna	dialects
dialog	dialogue
diamant	diamond
diamanter	diamonds
diameter	diameter
diamond	diamond
dianno	di'anno	dianno
dickens	dicken's
dickinson	dickinson
diego	diego
digerdöden	the black death
digital	digital
dikt	poem
diktator	dictator
diktatorn	the dictator	dictator
diktatur	dictator
diktaturen	dictatorship
dikter	poems
dillinger	dillinger
dimensioner	dimensions
din	your	yours
dinosaurier	dinosaurs
dinosaurierna	dinosaurs
diplomatiska	diplomatic
direkt	direct	directly
direkta	direct
direktör	director
diskar	disks
diskografi	discography
diskriminering	discrimination
diskussion	discussion
diskussioner	discussions
diskutera	discuss
diskuterades	discussed
diskuteras	discussed	is discucssed
diskuterats	been discussed	discussed
disney	disney
disneys	disneys	disney's
distinkt	distinct	distinctive
distinkta	distinct
distribution	distribution
distributioner	distributions
distrikt	district
distriktet	district
dit	there	where
ditt	your
dittills	thus far
diverse	some
division	division
divisionen	division
dj	dj
djup	deep
djupa	deep
djupare	depth	deeper
djupt	deeply	deep
djur	animals
djurarter	species of animals	animal species	species
djuren	the animals
djurens	the animals	animal
djuret	the animal
djurgården	djurgården
djurgårdens	djurgården's
djävulen	devil	the devil
dna	dna
dns	dns
dock	nevertheless	however
dog	died
doktor	doctor
dokument	files	documents
dokumenterade	documented
dokumentär	documentary
dollar	dollar
dom	judgement	conviction
domare	judge
domaren	the judge
domen	judgment	verdict; judgement
dominans	dominant	dominance
dominera	dominate
dominerade	dominated
dominerades	was dominated
dominerande	dominating
dominerar	dominates	dominate
domineras	dominated
dominerat	dominated
domkyrka	cathedral	abbey
domkyrkan	cathedral	the cathedral
domstol	court
domstolar	courts
domstolen	the court
don	don
donald	donald
donau	donau	the danube
donna	donna
dop	baptismal	baptism
dopamin	dopamine
dos	dosage
dotter	daughter
dottern	the daughter	daughter
downs	down
dr	doktor	dr	doctor
dra	pull; (with)draw
drabbade	suffering	affected
drabbades	affected	where hit by	afflicted
drabbar	affect	troubles	afflict
drabbas	suffer	troubled with
drabbat	affected
drabbats	affected	afflicted
drag	characteristic	move	trait; characteristic; feature
dragit	drawn	dragged
drama	drama
dramat	the drama
dramaten	dramaten
dramatiker	playwright	dramatist	dramatists
dramatiska	dramatic	dramatical
dramatiskt	dramatic	dramatically
dramer	dramas	plays
draperi	curtain	drapery; curtain	drapery	curtian
drar	earn	drag
dras	draw	make (assumptions, references)
dream	dream
drev	pursued	drove	led
drevs	concentrated	was driven
dricka	drink
dricker	drink	drinks
drift	drift
driva	operate	run
drivande	drive	driving
driver	driver	drive
drivs	driven	run
drog	draw	pulled
drogen	the drug	drug
droger	drugs
drogmissbruk	drug abuse, substance abuse, drug addiction	drug
drogs	was pulled	was
drottning	queen
drottningen	the queen
dryck	drinks
drycken	beverage	the drink
drycker	beverages
drygt	approximately
dräkt	costume	outfit
dröja	take
dröjde	was not until	not until
dröm	dream	syndrome
drömmar	dreams
dsmiv	dsm-iv
du	you
dubai	dubai
dubbel	double
dubbelt	double
dubbla	double
dublin	dublin
duett	duet
dvd	dvd
dvs	(det vill säga) namely that	i.e.
dvärg	dwarf
dvärgar	dwarves	dwarfs
dy	younger
dygn	day
dygnet	day
dyker	dives
dylan	dylan
dylikt	such
dynamiska	dynamic
dyrare	more expensive	expensive
dyraste	most expensive
dyrt	a high price	expensive	dearly
dä	the elder
däggdjur	mammalian	mammal
däggdjuren	the mammals
där	where	were
därav	thereof
därefter	then	thereafter
däremot	on the contrary	however, on the contrary	however
därför	because	therefore
däribland	among them	including
därifrån	from there
därigenom	by which	thereby
därmed	thus	consequently	therefore
därpå	darpa	thereon
därtill	thereto
därutöver	in addition	moreover
därvid	thus; thusly; then	therewith
då	then	when
dålig	poor
dåliga	bad
dåtidens	past times	yesterdays	that time
dåvarande	then	formerly
dö	die
död	dead	dod
döda	dead
dödad	killed
dödade	killed
dödades	killed	were killed
dödar	kills
dödas	killed
dödat	killed
döden	death
dödlig	lethal	mortal
dödligheten	mortality
dödligt	lethal	deadly
dödsfall	death
dödshjälp	euthanasy	euthanasia
dödsoffer	death victim	casualty	victim
dödsorsaken	cause of death
dödsstraff	death penalty
dödsstraffet	capital punishment; death penalty	the death penalty
dök	turned	dove
dömande	sentencing	judging
dömd	convicted	sentenced
dömdes	sentenced	was convicted
döpt	named	baptized
döpte	renamed
döptes	baptised	renamed	renamed; named
dör	dies	die
dött	died
döttrar	daughters
e	e
earl	earl
earth	earth
ebba	ebba
economic	economic	ecomomic
ecuador	ecuador
ed	ed
eddie	eddie
edgar	edgar
edison	edison
edith	edith
edmund	edmund
edvard	edvard	edward
edwall	edwall
edward	edward
edwards	edward's
edwin	edwin
effekt	effect
effekten	the effect	effect
effekter	effects; repercussions
effekterna	the effects	effects
effektiv	effective
effektiva	effective
effektivt	effective
efter	after
efterfrågan	demand
efterföljande	subsequent
efterföljare	following	follower
efterhand	hindsight
efterkrigstiden	the post-war period	post-war era
efternamn	last name	lastname
eftersom	while	because
efterträdare	successor
efterträddes	succeeded
eftervärlden	posterity	the world
efteråt	afterwards
egen	own
egendom	property
egenskap	trait	ability
egenskaper	characteristics	qualities
egenskaperna	the qualities	properties
egentlig	actual; factual; real	actual
egentliga	real one	actual
egentligen	really
eget	own
egna	own
egypten	egypt
egyptens	egypts	egypt's
egyptiska	egyptian
eiffeltornet	the eiffel tower
einstein	einstein
einsteins	einstein	once a	einsteins
ej	not	no
eker	united	spoker	spoke	spokes
eklund	eklund
ekman	ekman
ekologi	ecology
ekologiska	ecological
ekonomi	economic	economy
ekonomier	economies
ekonomin	the economy	economy
ekonomisk	economic
ekonomiska	economical
ekonomiskt	economic	economical
ekosystem	ecosystem	eco system
ekr	ad	ekr
ekvatorn	equator	the equator
eld	fire
elden	the fire
electric	electic
elektricitet	electricity
elektrisk	electric
elektriska	electrical
elektriskt	electric
elektromagnetisk	electromagnetic
elektron	electron
elektroner	electron	electrons
elektronik	electronics
element	elements
eleonora	eleonora
elever	students
eleverna	the pupils	the students
elin	elin
elisabeth	elisabeth
elit	elite
eliten	the elite
elitserien	elite series	elitserien
eller	or
elton	elton
elva	eleven
elvis	elvis
em	european championship
emellan	inbetween; between	between
emellanåt	once in a while	occasionally
emellertid	however
emi	emi
emigrerade	emigrated
emil	emil
eminem	eminem
emma	emma
emmanuel	emmanuel
emo	emo
empati	empathy
empire	empire
en	a
ena	one
enade	united
enades	agreed
enastående	exceptional
enat	united
enbart	only
encyclopedia	encyclopedia
enda	single	only
endast	only	merely
ende	only
energi	energy
energikälla	energy source	energy call
energikällor	energy resources	energy sources	sources of energy
energin	the energy	energy
energy	energy
engagemang	commitment
engagerad	dedicated	engaged
engagerade	dedicated	engaged	committed
engels	engels
engelsk	english
engelska	england	english
engelskan	the english	english
engelskans	english
engelske	the english	english
engelskspråkiga	english-speaking	the english language
engelsmännen	english people	the english	the british
england	england
englands	england's
english	english
enhet	unit	entity
enheten	the unit
enheter	units
enhetlig	unitary	uniform
enighet	unity
enkel	simple	plain
enkelt	easy
enkla	simple	single
enklare	easier	simpler
enklaste	the simplest	easiest
enlighet	according (to)	according
enligt	according (to)	according to
enorm	enormous
enorma	enormous
enormt	gigantic
ens	even	one's
ensam	alone
ensamma	alone
enskild	single
enskilda	individual
enskilt	individually
enstaka	occasional	single
entertainment	entertainment
enzymer	enzymes
ep	ep
epicentrum	epicentre
epok	epoch
epoken	the epoch
epost	e-mail	email
er	you	your
era	yours
eran	era
erbjuda	offer
erbjuder	offers
erbjöd	offered
erbjöds	offered
erektion	erection
erfarenhet	experience
erfarenheter	experiences	experience
erhållit	acquired	received
erhöll	obtained	recieved	acquire
eric	eric
ericsson	ericsson
erik	erik
eriksson	eriksson
eritrea	eritrea
erkänd	acknowledged
erkända	acknowledged	recognized
erkände	confession	acknowledged
erkänna	recognize
erkännande	recognition
erkänner	admits	recognize
erkänt	recognized
ernest	ernest
ernman	ernman
ernst	ernst
eros	eros
ersatt	replaced
ersatte	replaced
ersattes	was replaced by	replaced
ersatts	replaced	(has been) replaced
ersätta	replace
ersättare	replacement
ersättning	pay
ersätts	replaced
erövra	conquer
erövrade	conquered
erövrades	conquered	(was) conquered	concoured
erövring	conquest
erövringar	conquests
erövringen	conquest
estetik	esthetics
estetiska	aesthetic
estland	estland	estonia
estniska	estonian
et	et
etablera	establish
etablerad	established
etablerade	established
etablerades	established	was established
etablerat	established
etanol	ethanol
etik	ethics
etiken	the ethic	ethics
etiopien	ethiopia	ethiopian
etiopiska	ethiopian	etiopian
etiska	ehtical	codes
etnicitet	ethnicity	ethnic
etnisk	ethnic
etniska	ethnic
etniskt	ethnical
ett	a	one; a; an
etta	number one	first
etymologi	etymology
eu	eu
euro	euro
euron	the euro	euro
euroområdet	eurozone	convergence report
europa	europe
europacupen	euro (-pean) cup	european cup
europaparlamentet	european-parliament	the european parliament
europarådet	council of europe	european council
europas	europe
europe	europe
european	european
europeisk	european
europeiska	european
européer	europeans
européerna	europeans
eurovision	eurovision
eus	eu
eva	eva
evangelierna	the gospels
evangeliska	evangelical
evans	evans
evenemang	event
eventuell	any
eventuella	any	eventual
eventuellt	eventually	possibly
evert	everted	evert
everton	everton
eviga	eternal
evigt	forever	eternal
evolution	evolution
evolutionen	the evolution
evolutionsteorin	theory of evolution
ex	eg
exakt	accurately
exakta	exact
examen	exam
exempel	example	for example; for instance; sample(-s)
exempelvis	e.g.
exemplar	example	copies
exemplet	the example	example
exil	exile
existens	existence
existensen	existence
existera	exist
existerade	existed	existing
existerande	existing
existerar	exists
existerat	existed
exklusiv	exclusive
expandera	expand
expansion	expansion
expansionen	the expansion
expedition	expidition	expedition
expeditionen	the expidition	expedition
expeditioner	expeditions
experiment	experiment
experimenterade	experimented
experter	experts
explosionen	the explosion
export	export
exporten	exports	the export
express	express
expressen	expressen
externa	external
extra	optional
extrem	extreme
extrema	extreme
extremt	extreme
fabriker	factories
facebook	facebook
fackföreningar	unions
facto	facto
facupen	fa cup	fa-cup
fader	father
fadern	the father
faderns	the father's
fagocyt	phage	fagocyte	phagocyte
fakta	fact
faktiska	actual
faktiskt	in fact; actually; indeed	actually	really
faktor	factor
faktorer	factors
faktorn	factor
faktum	fact
fall	where
falla	fall
fallen	cases
faller	fall
fallet	the case
fallit	fallen
falska	false
falskt	false
familj	family
familjen	the family
familjens	the familys
familjer	families
familjerna	families
fan	devil
fann	found
fanns	was
fans	fans
fansen	fans
far	father
fara	danger
farbror	uncle
farfar	paternal grandfather
farlig	dangerous	hazardous
farliga	dangerous
farligt	dangerous
fars	father's	father
fart	speed
fartyg	ship; vessel	ship
fartyget	ship; vessel
fas	phase
fascism	fascism
fascismen	the fascism	fascism
fascisterna	fascists
fascistiska	fascist	fascistic
fasen	phase
faser	phase	phases
fast	though; although; fixed; permanent	even though
fasta	firm; set; solid; fast; fasting
fastigheter	real estates
fastlandet	mainland
fastställa	determine	confirm
fastställdes	confirmed
fastän	although
fat	fat
fatta	make
fattas	taken
fattiga	poor
fattigare	poorer
fattigaste	the poorest	poorest
fattigdom	poverty
fattigdomen	poverty
fauna	fauna
fbi	fbi
fc	fc
fci	fci
fd	ex
feber	fever
februari	februari	february
federal	federal
federala	federal
federation	federation
federationen	federation	the federation
fel	faults	errors	error
felaktig	incorrect	false
felaktiga	false
felaktigt	incorrect	erronenous
felix	felix
fem	five
feminism	feminism
feminismen	feminism
feminister	feminists
feministiska	feminist
femte	fifth
femton	fifteen
fenomen	phenomenon	phenomenazaqq
fenomenet	the phenomenon	phenomenon
feodala	feudal
ferdinand	ferdinand
fermentering	fermentation
fernando	fernando
fest	party	fest
fester	parties
festival	festival
festivalen	festival	the festival
festivaler	festivals
fett	fat
ff	ff
fick	got	was
fiende	enemy
fienden	enemy	the enemy
fiender	enemies
fifa	fifa
figur	figure
figuren	the character	figure
figurer	figures
figurerna	figures	characters
fiktion	fiction
fiktiv	fictive
fiktiva	romantic
fil	master of
filip	phillipe	filip
filippinerna	the philippines
film	film
filmatiserats	cinematized	screened
filmen	the movie	film
filmens	the film's	film
filmer	films	movies
filmerna	the movies
filmografi	filmography
filosofen	the philosopher
filosofer	philosophers	philosopher
filosofi	philosophy
filosofin	philosophy	the philosophy
filosofins	philosophy	the philosophy
filosofisk	philosophic
filosofiska	philosophical
fina	beautiful	fine
final	final	finite, final
finalen	final
finansiella	financial
finansiera	fund	finance
finansieras	financed	finansed
finansiering	financiation
finanskrisen	financial crisis	the financial crisis
finger	finger
fingrar	fingers	finger
finland	finland
finlands	finlands
finländska	finish	finnish
finna	found
finnas	found	(be) found	exists
finner	finds
finns	exist	there is
finsk	finnish
finska	finnish
fira	celebrate
firade	celebrated
firades	was celebrated
firandet	celebrate	the celebration
firar	celebrates	celebrate
firas	celebrated	celebrate
fire	fire
fisk	fish
fiskar	fishes
fiske	fishing
fission	fission
fjorton	fourteen
fjädrar	feathers
fjärde	fourth
fjärdedel	quarter	fourth
flagga	flag
flaggan	the flag
flaggor	flags
flames	flames
flamländska	flemish
flandern	flanders
fler	more
flera	many	multiple
flertal	several	majority group
flertalet	majority; plurality	several
flest	most	the most
flesta	most
flicka	girl
flickan	girl	the girl
flickor	girls
flickvän	girlfriend
flight	flight
flitigt	actively	frequent
flod	river
floden	the river
floder	rivers
floderna	floods	the rivers
flora	flora
florens	florence	florens
florida	florida
flotta	fleet
flottan	the fleet	navy	the navy
floyd	floyd
fly	escape
flydde	fled
flyg	airforce
flyga	fly
flygande	flying
flygbolag	airline
flyger	flies	flying
flygplan	airplane
flygplats	airport
flygplatsen	the airport
flygplatser	airports	air ports
flygvapnet	air force	the airforce
flykt	escape
flyktingar	refugees
flyr	flees	escapes
flytande	floating	liquid
flyter	flows
flytt	escaped	fled
flytta	move
flyttades	moved
flyttar	move
flyttas	is moved	moved
flyttat	moved
flöde	feed
flög	flew
fn	un	the un
fns	un's	tris
fokus	focus
fokusera	focus
fokuserade	focused
fokuserar	focuses	focus
folk	public	people
folke	folke
folken	the peoples
folket	the people
folkets	the people's
folkgrupper	ethnic groups
folklig	popular
folkliga	popular	folk
folkmord	genocide
folkmordet	genocide
folkmun	popular lore; popularly	colloquially	common speech
folkmusik	folk music
folkmängd	population size	population
folkmängden	population
folkomröstning	referendum
folkpartiet	peoples party
folkrepubliken	people's republic	people"s republic
folkrikaste	populous	people rich	most populus
folkräkning	head count
folkräkningen	census
folkslag	kind of people	peoples
folktro	popular belief	folklore
folkvalda	elected	popularly elected
fontsizes	fontsizes
football	football
force	force
ford	ford
fordon	vehicle/-s	vehicles	vehicle
form	form
format	format	shaped
formatet	the format	size	format
formel	formula
formell	formal
formella	formal
formellt	formally
formen	the form
former	forms
formerna	forms
forna	former
fornnordiska	old nordic	ancient nordic
forntida	pristine	prehistoric
forsberg	forsberg
forskare	researcher	researchers	scientists
forskaren	researcher
forskarna	the scientists	scientists
forskning	research
forskningen	the science
fort	quickly
fortfarande	still
fortplantning	reproduction
fortsatt	further	continued
fortsatta	continued
fortsatte	continued
fortsätta	remain	continue
fortsätter	continues	continue
fortsättning	continuation
fortsättningen	the continuation
forum	forum
fossil	fossil
fossila	fossilized	fossil
foster	embryo	fetus	fetuses	foster	embryonic	fetal
fot	foot
fotbeklädnad	chaussure	foot gear	shoewear	chausurre	footwear
fotboll	football
fotbollen	soccer	football
fotbollslandslag	football team	national football team
fotbollsspelare	football player	footballers
foten	foot
fotnoter	footnotes
foto	photo
fotografier	photographs
foton	photos
fotosyntesen	photosynthesis
fragment	fragment
fralagen	the fra law
fram	until	out
framför	in front of	above
framföra	express	convey
framförallt	in particular; above all	above all
framförde	performed	presented
framfördes	framfordes
framförs	is presented	performed
framfört	expressed	presented
framförts	forward	performed
framgång	success
framgångar	successes	success
framgångarna	the successes
framgången	the success
framgångsrik	successful
framgångsrika	successful	succesful
framgångsrikt	successful	successfully
framgår	will be seen	clear	is shown
framsteg	progress
framställa	represent; depict; produce	the installation
framställning	production
framställs	is depicted	prepared
framstående	prominent
framtid	future
framtida	future
framtiden	future	the future
framträdande	apperance	appearance
framträdanden	appearances
framträdde	appeared
framträder	stand	appear
framåt	forward	forth
francis	francis
francisco	fransisco
franco	franco
franklin	franklin
frankrike	france
frankrikes	frances	france's
fransk	french
franska	french
franske	the french	french
franskt	french
fransmännen	the french	french
franz	franz
français	francais
fred	peace
freddie	freddie
freddy	freddy
freden	the peace	peace
fredliga	peaceful
fredrik	fredrik
fredsbevarande	peacekeeping
fredspris	peace prize
fredspriset	peace prize	peace price	nobel peace prize
freedom	freedom	frihet
freja	freja
frekvens	frequencies	frequency
freud	freud
fri	free
fria	free
friedrich	friedrich
frigörelse	liberation
frigörs	released	is released
frihet	freedom
friheten	freedom; liberty	liberty
frihetliga	libertarian
friidrott	track and field
frisk	healthy	fresh
friska	healthy	fresh	healty
fristående	independent	stand-alone
fritid	free time	recreational	leisure	leisure time	freetime	spare time	leisure time; spare time
fritt	free
fritz	fritz
frivillig	optional
frivilliga	volunteers	optional
frivilligt	voluntarily	voluntary
frodo	frodo
from	from
front	front
fronten	front	the front
fru	mrs.	wife
frukt	fruit	fruits
fruktade	feared
frälsning	salvation
främja	further	promote
främmande	foreign; alien	undesirable	foreign
främre	front
främst	foremost; primarily; chiefly	primarily
främsta	primary; foremost; primarily; principally	request
främste	chief	premier
fråga	fraga	ask	question
frågade	asked
frågan	the question
frågor	questions
frågorna	questions; issues
från	from
frånträde	relinquishment	withdrawal
frånvaro	absent	absence
fröken	miss
fröväxter	seed-bearing plants	seed plants	phanerogams	seed plant	spermatophytes	spermatophyte
fss	fss
fuglesang	fuglesang
fuktiga	damply
fuktigt	moist	humid
full	full
fulla	full	complete
fullständig	full	complete
fullständiga	complete
fullständigt	completely	full
fullt	full; fully; completely	completely	full
fungera	act
fungerade	working
fungerande	functioning	effective	working
fungerar	functions	works
funktion	function
funktionella	functional
funktionen	function	the function
funktioner	functions
funktionerna	functions	the functions
funnit	found
funnits	been
fursten	prince
fusion	fusion
fusionen	the fusion
futharkens	futhark	the futhark's
fylla	fill
fyllde	completed	filled
fyller	turns	turn; fill
fynd	finding; finds
fynden	finds; findings	findings
fyra	four
fyrtio	forty
fysik	physics
fysikaliska	physical
fysiker	physicist
fysiologi	physiology
fysiologiska	physiological
fysisk	physical
fysiska	physical
fysiskt	physically	physical
fält	field
fältet	the field	field
fälttåg	crusade	campaign
fängelse	prison
fängelsestraff	imprisonment	prison
fängelset	prison
fängslade	inprisoned	confine	imprisoned
fängslades	imprisoned; jailed, gaoled; incarcerated	jailed
färdas	travels
färdig	done
färdiga	completed
färg	colour	colors
färgade	colored
färgen	the color
färger	colors
färgerna	colors
färre	less
färöarna	faroe islands	the faroe islands
fäste	bracket	attachment
fästning	fortress
få	have; make; few	fa
fåfotingar	fafotingar	pauropoda	pauropods
fågel	bird
fågelarter	species of bird
fågelhundar	bird dogs
fåglar	birds
fåglarna	the birds	birds
fåglarnas	the birds'	birds
fånga	capture
fångar	prisoners
fångenskap	captivity
får	can	allow
fåtal	a few
fått	was given	with
föda	give birth; food	give birth
född	born
födda	born
födde	gave birth too	born
föddes	was born	born
födelse	birth
födelsedag	birthday
födelsetal	birthrate	birth rate
föder	give birth of	gives birth
föds	born
födseln	birth	the birth
föga	little	hardly; little
följa	following	follow
följaktligen	consequently
följande	following	the following
följas	followed
följd	effect
följde	followed
följden	result	the cause
följder	impact	consequences
följdes	followed	was followed
följer	resulting
följeslagare	companion
följs	followed
följt	followed
föll	fell
fönster	windows	window
för	of	to; for	for
föra	pre	lead
föranledde	brought about	led
föras	be	be brought	taken to
förband	units; formations; bound (themselves)	bond
förbi	past	past the	pass
förbindelse	connections	connection
förbindelser	connections	relations
förbinder	connects	undertake
förbjuda	ban	forbid
förbjuden	smoking
förbjuder	prohibiting	forbids
förbjudet	prohibited
förbjudna	forbidden	prohibited
förbjöd	forbid
förbjöds	forbidden
förblev	remained
förblir	remains	remain
förbränning	combustion
förbud	ban	prohibition
förbudet	ban	the union
förbund	union	league; alliance; union; compact; covenant
förbundet	the union
förbundskapten	manager
förbundsrepubliken	the federal republic	federal republic
förbundsstat	federal state
förbättra	improve
förbättrade	improved
förbättringar	improvements	improvement
förde	led
fördel	advantageously	advantage
fördelade	divided	distributed
fördelar	advantages	share
fördelas	distribute	distributed
fördelen	advantage	the advantage
fördelning	distribution
fördelningen	distribution
fördes	sea were entered
fördomar	bias	prejudice	prejudices
fördrag	agreement	treaty
fördragen	treaties	the compacts
fördraget	the treaty	treaty
fördrevs	was banished	ford described	driven away
före	ahead (of), before
förebild	role model
förebyggande	preventing	preventive
föredrar	prefer
föredrog	prefered	preferred
förefaller	appear
föregående	preceeding; previous	previous
föregångare	predecessor
föregångaren	predecessor
förekom	was
förekomma	occur	be found
förekommande	occuring
förekommer	preferred is	occurs
förekommit	occured	occurred
förekomst	presence
förekomsten	existence	presence
föreligger	is	exist
föremål	object	subject
förena	combine	unite
förenade	united
förening	union
föreningar	associations	organizations
föreningen	association	the association
förenklat	simplified	made easier
förenta	united
föreslagit	suggested	proposed
föreslagits	was suggested
föreslog	suggested	propose
föreslogs	was suggested
föreslår	suggest
förespråkade	advocate	advocated
förespråkar	advocate
förespråkare	spokesman
föreställa	imagine	pretend; imagine
föreställande	depicting
föreställer	picture	depicts
föreställning	performance
föreställningar	performances	notions
föreställningen	the idea	the concept	show
företag	company	companies
företagen	the companies
företaget	the company
företagets	the company's	the corporation's
företeelse	experience; phenomenon; feature	phenomenon
företeelser	phenomena
företrädare	representatives
företräder	preferred trades	representing
författare	author
författaren	the author
författarna	the authors	writers
författarskap	the writer	authorship
författning	constitution
författningen	constitution
förfäder	ancestors
förföljelse	persecution
förföljelser	pursuits	persecutions
förgäves	in vain
förhandla	negotiate
förhandlingar	negotiations
förhandlingarna	the negotiations	negotiations
förhindra	prevent
förhindrar	prevents
förhistoria	prehistory
förhistorisk	forhistorisk	prehistorian
förhärskande	dominant	prevailing
förhållande	in relation	(in) comparison (to)
förhållanden	relationships	conditions
förhållandena	conditions	the conditions
förhållandet	the ratio	relationship
förhållandevis	relatively
förhåller	relate	relates
förhöjd	enhanced
förintelsen	the genocide
förklara	explain
förklarade	explained	said
förklarades	was explained
förklaras	explained
förklarat	declare
förklaring	explaination	explanation
förklaringar	explanations
förklaringen	the explanation
förknippad	associated
förknippade	associated
förknippas	associated to	associate
förkortas	abbreviated
förkortat	shortened
förkortning	abbreviation
förkortningar	abbreviations
förlag	magazine
förlaget	publisher	the publisher
förlopp	process	pattern	developments
förlora	lose
förlorade	lost
förlorades	was lost
förlorar	loss	loses
förlorat	lost
förlust	loss
förlusten	loss	loss; defeat
förluster	losses
förlusterna	the losses
förlängning	overtime; extension; prolongation	extension
förlängningen	elongation
förmedla	pass; express; mediate	pass
förmodligen	probably	presumably
förmåga	abilities	ability
förmågan	the ability
förmågor	capacities	abilities
förmån	benefit	advantage; in favor of; benefit
förmögenhet	fortune	wealth
förnuft	reason
förnuftet	reason	the common sense
förorter	suburbs
förr	sooner; past	sooner	before
förra	last	former
förrän	until	before
förs	led	rapids
församling	congregation
församlingar	parishs	assemblies
församlingen	parish	congregation
förslag	proposal	'proposal
förslaget	proposition	the suggestion
först	first
första	first
förstaplatsen	first place
förste	chief	the first
förstnämnda	first-named	aforementioned	first named
förstod	understood
förstärka	strengthen
förstå	understand	first
förståelse	understanding
förståelsen	the understanding
förstår	understand	forstar
förstås	course	mean:
förstöra	destroy	ruin; destroy
förstördes	was destroyed
förstörelse	destruction
försvann	disappeared
försvar	defence
försvara	defend
försvarade	defended
försvarare	defender
försvaret	repository	the defense
försvarets	defense	forsvarets	the defence's
försvarsmakt	armed forces
försvarsmakten	national defence	national defense
försvarsminister	minister of defence
försvinna	vanish	disappear
försvinner	disappears	disappearing	disappear
försvunnit	disappeared
försäkra	make sure	insure
försäljning	sale	sales
försäljningen	sales
försämrades	worsened	worsening
försök	expirements
försöka	try	attempt
försöken	attempts	the tries
försöker	try	tries	trying
försökt	tried
försökte	try	tried
försörja	support
försörjde	provided
försörjning	sustention	sustentation
fört	led	lead
förteckning	index	listing	label
förtjust	fond	delighted
förtroende	confidence	trust
förtryck	opression
förts	brought	cont
förut	before
förutom	besides; in addition to; aside from
förutsätter	assume	assumes
förutsättning	prerequisite
förutsättningar	prerequisites	(pre-)conditions	condition
förutsättningarna	prerequisites
förvaltning	management	administration
förvaras	is stored
förväntade	expected
förväntas	expected
förväntningar	expectations
förväxla	mistake
förväxlas	mixed up (with)	confused	mistaken
föräldrar	parents
föräldrarna	the parents
förälskad	in love
förändra	change; alter; replace	change
förändrade	changed
förändrades	changed
förändras	changes
förändrats	changed
förändring	change
förändringar	changes
förändringarna	changes	change
förändringen	the change
förödande	devastating
fötter	feet	on its feet
fötterna	feet	the feet
fötts	born	borned
führer	fuhrer	fuehrer
gabriel	gabriel
gaga	gaga
galax	galaxy
galaxer	galaxies
galilei	galilei
galileo	galileo
gallagher	gallagher
galleri	gallery
gallien	gaul
gamla	ancient	old
gamle	old
gammal	old
gammalt	old
gandalf	gandalf
gandhi	gandhi
gandhis	gandhi's
ganska	fairly	quite
garantera	guarantee
garanterar	ensures
garvey	garvey
gary	gary
gas	gas
gasen	gas
gata	street
gatan	the street
gates	gates
gator	streets
gatorna	the streets
gav	gave
gavs	gave
gaza	gaza
gazaremsan	gaza strip	the gaza strip
ge	to give	give
gemensam	joint	common
gemensamma	joint	common
gemensamt	in common
gemenskap	fellowship
gemenskapen	the collective	community
gemenskaperna	communities	community
gen	gene
genast	immediately	at once
genen	gene	the gene
gener	genes
general	general
generalen	the general
generalguvernören	governor-general	governor general	general governor
generalsekreterare	the secretary-general	secretary general
generation	generation
generationen	generation	the generation
generationer	generations
generell	general
generella	overall	general
generellt	generally
generna	genes	the genes
genetik	genetics
genetisk	genetic
genetiska	genetic
genetiskt	genetically	genetic
genom	through
genombrott	breakthrough
genombrottet	break-through	breakthrough
genomför	implement	carry out
genomföra	perform	out
genomföras	be performed	carry out
genomförde	carried out
genomfördes	was	was carried out
genomförs	implemented, carried through	conducted
genomfört	carried out	implemented	carried through
genomförts	out
genomgick	underwent
genomgripande	good	comprehensive; radical
genomgående	consistently	pervading
genomgår	undergoes	undergoing
genomgått	experienced	passed
genomslag	breakthrough
genomsnitt	average
genomsnittet	average	the average
genomsnittlig	average
genomsnittliga	average
genre	genre
genren	genre
genrer	genres
gentemot	towards	against
genus	gender	genus
geografi	geography
geografisk	geographic	geographical
geografiska	geographical	spatial
geografiskt	geographically	geographic
geologi	geology
geologiska	geological
geologiskt	geological
geomorfologi	geomorphology
georg	georg
george	george
georges	georges
georgien	georgia
georgier	the georgians	georgian	georgians	georgier
ger	gives; is giving	give
germanska	germanic	germanian
ges	given	be given
gestalt	character	figure
gestalter	beings	figures
gett	given	gave
ghana	ghana
gia	gia
gick	went	passed
gift	married
gifta	marry	married
gifte	married
gifter	marries
giftermål	marriage	marrige
giftsnokar	elapidae	venomous conks	venomous grass snake	venomous snakes	elapidaes	poisonous snakes	venomous snake	elapids	venom snooping
gigantiska	gigantic
gillade	liked	approved; liked
gillar	likes	enjoy; like
giovanni	giovanni
girl	girl
girls	girls
gisslan	hostage
gitarr	guitar	guitarr
gitarrist	guitarist
gitarristen	the guitarist
givaren	donor	the giver	dealer
given	given
givet	granted
givetvis	naturally
givit	gave
givits	given
gjord	made
gjorda	made	done
gjorde	did
gjordes	made	was made
gjort	made	created
gjorts	done
glad	happy
glada	happy
glas	glass
glenn	glenn
global	global
globala	global
globalt	globally
globe	globe
globen	the globe
gloria	gloria
glukos	glucose
glädje	joy
glödlampor	lightbulbs	light bulbs
go	go
god	good
goda	good
godkände	approved
godkändes	approved
godkänna	approve
godkännande	approval	authorization
godkännas	pass on	approved	be approved
godkänt	approved
gods	domain	goods
goebbels	geobbels
gogh	gogh
golf	golf
golvet	the floor
gom	palate	mouth	roof of mouth	gum
google	google
gorbatjov	gorbachev	gotbatjov
gordon	gordon
got	got
gotiska	gothic
gotland	gotland
gotlands	gotland's
gott	practically; good
grace	grace
grad	grade	rate
graden	rate	the degree
grader	degrees
gradvis	gradually
grafit	graphite
graham	graham
grammatik	grammar
grammis	grammy
grammy	grammy
gran	spruce
grand	grand
grande	grand
grannar	neighbours
granne	neighbour	neighbor
grannlandet	the neighbouring country
grannländer	neighboring countries	neighboring lander
grannländerna	neighbors	neighbouring countries
granska	review
granskning	review
grant	word
gratis	free
grav	grave
graven	the grave	grave
gravid	pregnant
graviditet	pregnancy
graviditeten	the pregnacy	the pregnancy
gravitation	gravitation
gray	gray
greker	greek	greeks
grekerna	greeks	greek
grekisk	greek
grekiska	greek
grekiskans	the greek's	greek
grekland	greece
greklands	greece's
gren	branch
grenar	branches
grenen	the branch	branch
greps	was arrested	(was) arrested
greve	earl
griffin	griffin
griffon	griffon
grovt	heavy	roughly
grund	in the context: "på grund" = because of	because
grunda	found	base
grundad	founded
grundade	founded	based
grundades	founded	was founded
grundande	founding
grundandet	founding (of)	founding
grundar	bases
grundare	founder
grundaren	the founder	founder
grundarna	founders
grundas	is based	based
grundat	founded	(was) found	based
grunden	base
grunder	bases
grundlag	constitution
grundlagen	constitution	the constitutional law
grundläggande	primary	fundamental
grundskolan	elementary school
grundämne	element
grundämnen	elements
grundämnet	the element	element
grupp	group
gruppen	the group
gruppens	group (-s)	group
grupper	groups
grupperingar	groups	groupings
grupperna	groups
gruppspelet	groupplay	group play
gräns	limit	border
gränsar	border	borders (to)
gränsen	border
gränser	borders
gränserna	borders	the borders
gräs	grass
gräslök	chive	chives
grå	gray	grey
grön	green
gröna	green
grönland	greenland
grönsaker	vegetables
grönt	green
grönwall	grönwall
guatemala	guatemala
gud	god
gudar	gods
gudarna	the gods
gudarnas	the gods'	god's
guden	the god
gudinnan	the godess
gudom	deity
gudomlig	divine
gudomliga	divine
guds	god's
guevara	guevara
guide	guide
guillou	guillou
guinea	guinea
gul	yellow
gula	yellow
guld	gold
guldbollen	golden ball	guldbollen
gunnar	gunnar
guns	guns
gunwer	gunwer
gustaf	gustaf
gustafs	gustafs	gustaf's
gustafsson	gustafsson
gustav	gustav
gustavs	gustavs	gustav
guvernör	governor
guyana	guyana (name)	guyana
gyllene	golden	golden; gilded
gymnasiet	high school	gymnasium
gymnasium	high school
gälla	be valid
gällande	regarding
gällde	applied	applied to
gäller	of	refer to	grating
gäng	group
gänget	the group	the gang
gärna	i'd love to	readily
gärning	deed
gärningar	deeds
gärningsmannen	perpetrator; offender	the offender	culprit
gäst	guest
gäster	guests
gävle	gävle
gå	go
gång	time	once
gången	time
gånger	times
gångna	past	past; gone
går	is	goes
gård	farm	house
gården	courtyard; house; farm (-house)
gått	gone	passed
gåva	gift
gör	does	makes
göra	do	do; doing
göran	göran	request
göras	made	be made	be made through
göring	goring
görs	made	is made to
gösta	gösta
göta	göta
götaland	götaland	gotaland
göteborg	gothenburg
göteborgs	gothenburg	gothenburgs
h	h
ha	be	have
haag	haag	the hague
haber	haber
haddock	haddock
hade	had
haft	had
haile	haile
haiti	haiti
hall	hall
halland	halland
halloween	halloween
hallucinationer	hallucinations
halmstad	halmstad's
halmstads	straw city	halmstad's
hals	throat
halsen	the throat
halt	stop; level	stop
halv	half
halva	half
halvan	the half
halvklotet	hemisphere
halvt	half
halvön	the peninsula
hamas	hamas
hamburg	hamburger
hamilton	hamilton
hamlet	hamlet
hammarby	hammarby
hamn	harbor	harbour
hamna	end
hamnade	landed	ended up
hamnar	lands	ports
hamnat	got	ended up	got in to
hamnen	harbour	the harbour
hampa	hemp
han	he
hanar	males
hand	care	hand
handboll	handball
handel	trade
handeln	trade; commerce	trade
handels	trade
handelsmän	merchants
handelspartner	trading partner
handen	the hand	hand
handla	act; buy; consume
handlade	was (about); traded
handlande	action
handlar	is	concerns
handling	act
handlingar	actions
handlingen	hand-writing	the plot	the story
hanen	the cock	the male
hanhon	he/she
hann	reached	managed to (in a period of time)
hannah	hannah
hannar	males
hans	his
hansson	hansson
hantera	handle
hantverk	crafting
hantverkare	handy worker	craftsman
har	is	has	have
harald	harald
harris	harris
harrison	harrison
harry	harry
hasch	hashish
hastighet	speed
hastigt	rapidly	fast
hat	hatred
hatar	hate	hates
hav	seas	sea	ocean
have	have
haven	the seas
havet	sea
havets	the seas
havs	at sea
havskattfiskar	catfishes	goatfish	catfish fish	catfish fishing	catfished	catfish	wolffish	have duty fish	mullet	seawolf	sea wolfs
havsnivån	sea level
hawaii	hawaii
hawking	hawking
hc	h.c.	h.c
hdmi	hdmi
he	he
heart	heart
heath	heath
heaven	heaven
hebreiska	hebrew
hedersdoktor	honorary doctor	honorary degree
hegel	hegel
heinrich	heinrich
heinz	heinz
hel	(whole) lot (of)
hela	entire
helena	helena
helgdagar	holidays
helhet	entirety	whole
helig	holy
heliga	holy	holy; holy
helige	holy
heligt	holy
helium	helium
hell	hell
heller	neither; nor
hellre	rather
hells	hells
hellström	hellström	hellstrom
helsingborg	helsingborg
helsingborgs	helsingborg's
helsingfors	helsingfors	helsinki
helsingör	helsingor	helsingör
helst	anyone	rather
helt	totally
helvetet	the hell
hem	home
hemingway	hemingway
hemland	homeland
hemlandet	the home country	the homeland
hemlig	secret
hemliga	secret
hemlighet	secretly
hemligt	secret
hemma	home	at home
hemmaarena	home ground
hemmaplan	home	home turf; domestic (level)
hemmet	the home
hemsida	homepage
hendrix	hendrix
henne	she	her
hennes	her
henri	henri - it's a name	henri
henrik	henrik
henriks	henry
henry	henry
hepatit	hepatite	heptatitis
herbert	herbert
hercegovina	herzegovina
hergé	herge	hergé
heritage	heritage
herman	herman
hermann	hermann
heroin	heroin	heroine
herr	mister	mr
herrar	gentlemen	men
herre	lord	master; lord
herren	the lord
herrens	lord
herrlandskamper	men's international contest	men's international contests
herrlandslag	men's national team
hertig	duke
het	hot	up to date
heta	hot	be named; be called	be called
heter	(is the) name (of)	is named
hett	hot
hette	named
hexadecimalt	hexa-decimal	hex
heydrich	heydrich
high	high
himlakroppar	celestial bodies
himlen	heaven
himmel	heaven
himmler	himmler
himmlers	himmlers
hinder	obstacle	barrier
hindra	hinder	prevent
hindrade	prevented	preventing
hindrar	prevents	stop; prevent
hindu	hindu
hinduer	hindu
hinduiska	hindu
hinduism	hinduism
hinduismen	hinduism
hinner	reach it (in time)	have time to
hiroshima	hiroshima
his	his
hisingen	hisingen
historia	history
historien	history
historiens	historys
historier	stories	history
historik	history
historiker	historians
historikern	historian
historisk	historic	historical
historiska	historical
historiskt	historic	historically	historical
history	history
hit	to here	here
hitler	hitler
hitlers	hitlers
hits	hits
hitta	see	make up	come up, find
hittade	found
hittades	was found
hittar	finds
hittas	found
hittat	found
hittats	found
hittills	date	so far
hiv	hiv
hjalmar	hjalmar
hjälp	help
hjälpa	helping
hjälper	helps	shows
hjälpmedel	aid	resources
hjälpt	helped
hjälpte	helped
hjärna	brain
hjärnan	brain	the brain
hjärnans	brain
hjärta	heart
hjärtat	heart	the heart
hms	hms
ho	ho
hockey	ice hockey	hockey
holland	holland
hollywood	hollywood
holländska	dutch
holm	holm
homo	homo	gay
homogen	homogenous
homosexualitet	homosexuality
homosexuell	homosexual
homosexuella	homosexual	gay
hon	she
honan	the female	female
honom	his	him
honor	ära
hopp	hopes	hope
hoppa	skip	drop out
hoppade	jumped
hoppades	hoped
hoppas	hope
hormoner	hormons
horn	horn	horns
hos	in; with	with
hotad	threatened
hotade	threatened
hotar	threatens
hotel	hotel
hotell	hotel
hotellet	the hotel
hotet	the threat	the threath
house	house
houston	houston
hov	court
hovet	court	the court
hovrätten	the court of appeal
how	how
howard	howard
hud	skin
huden	skin
hudfärg	color
hughes	hughes
hugo	hugo
human	human
humanism	humanistic	humanism
humanismen	humanism
humanistiska	humane	humanistic	humanist
humle	hop
humor	humour
humör	temper	mood
hund	dog
hundar	dogs
hunden	the dog	dog
hundra	hundred	one hundred
hundraser	alternative strains	breed of dogs
hundratal	hundred
hundratals	hundreds of	hundreds
hundratusentals	hundreds of thousands
hunnit	reached	had time to
hur	how	cage
huruvida	whether
hus	house	housing	a house
husen	housing	the houses
huset	the house
hushåll	household
huskvarna	huskvarna
hussein	hussein
hustru	wife
hustrun	the wife	his wife
huvud	head	main
huvudartikel	main article	principal article
huvuddelen	main part
huvudet	head	the head
huvudkontor	central office	headquarters
huvudort	main town	principal town
huvudperson	main person; main character	main character
huvudrollen	the main role	leading part
huvudsak	in principal; chiefly	main thing
huvudsakliga	main
huvudsakligen	generally	primarily
huvudstad	capital city
huvudstaden	capital
huvudstäder	capital cities	capitals
huvudvärk	headache
huxley	huxley
hyllade	celebrated
hyllning	tribute; homage
hypotes	hypothesized	hypothesis
hypotesen	the hypothesis	hypothesis
hypoteser	hypotheses	hypothesis
hyser	has	accomodates	holds
häcklöpning	hurdles	hurdles race	hurdling	hurdle	hacklopning	hurdle race	hurdle-race
hälft	half
hälften	half
hällristning	petroglyph	stone carving	rock carving	rock engraving	chives	rock carvings	rock	rock engravings
hälsa	tell (him i said hi)
hämnd	revenge
hämta	retrieve	fetch
hämtade	brought
hämtar	download	is	gets
hämtat	collected	taken
hända	may
hände	happened
händelse	event
händelsehorisonten	event horizon	the event horizon
händelsen	the occurence	event
händelser	handelsar	happenings
händelserna	the events	the happenings
händer	happens	hands
händerna	hands
hänga	hang
hänger	depends	hanger
hänsyn	consideration
hänt	suspension	happened
hänvisa	refer
hänvisade	refer
hänvisar	reference
hänvisning	reference
här	this; here	here
härifrån	from here	here
härkomst	origin
härledas	derived
härrör	derived
härskare	ruler
härstamma	originate	stem
härstammar	derived	stems
härstamning	origin	descent
häst	horse
hästar	horses
hästen	the horse
hästens	horses	horse's
hävda	claim
hävdade	claimed
hävdar	assert	maintain
hävdat	claimed
håkan	chin
håkansson	hakansson
hål	hole	hal
hålet	hole; gap	the hole
håll	ways	hold
hålla	keep
hållas	be held
håller	holds
hållet	way
hållit	held	maintained	kept
hållning	position	attitude
hålls	maintaned	is held
hår	hair
hård	diffcult	hard
hårda	hard
hårdare	harder	tougher
hårdast	the most	the hardest
hårdrock	hard rock
hårdrocken	hard rock
hårdvara	hardware	hardwere
håret	the hair
hårt	hard	resin
höftledsgrop	acetabulum	aetabulum	hip pit	hip joint fossa	hoftledsgrop
hög	high
höga	high
höger	right
högkvarter	headquarters	head quarter
höglandet	highlands	the highland
högra	right
högre	higher
högskola	college
högskolan	hogs school	university	college
högskolor	colleges
högst	highest	maximum
högsta	highest
högste	supreme	highest
högt	high	highly
högtid	festival	festival; holiday
högtider	holiday	feasts
högtryck	high pressure	pressure	anticyclone	high presssure
höja	hoja	increase	raise
höjd	height; above	height
höjder	altitudes	heights
höjdes	increased	was raised
höjdpunkt	highlight	climax	high point
höjer	rises	raising
höll	hold	gave
hölls	was held	was
hör	belong	hears
höra	hear
hörde	heard
hörn	corner
hörs	heard
hört	heard	heared
höst	autumn
hösten	the fall	the autumn
i	of	in
ian	ian
iberiska	iberian
ibland	sometimes
ibm	ibm
ibn	ibn
ibrahimović	ibrahimovic
icd	icd
icke	non	none
ida	ida
idag	today
ideal	ideals	ideal
identifiera	identification
identifierade	identified
identisk	identical
identitet	identity
ideologi	ideology
ideologier	ideologies
ideologin	the ideology
ideologiska	ideological
ideologiskt	ideologically	ideological
idol	idol
idrott	sports
idéer	ideas
idén	the idea	idea
ifall	if
ifk	ifk
ifråga	with regards to	in question
ifrågasatt	questioned
ifrågasatts	is questioned	questioned
ifrån	off
igelkott	hedgehog
igelkottar	hedgehogs
igelkotten	the hedgehog
igelkottens	the hedgehog's	hedgehog
igen	again	recognize
igenom	through
igång	start	start up
ihop	up	together
ihåg	remember
iii	iii
iiis	iii's	3's
iis	ii's
ikea	ikea
ikon	icon
illa	bad
illegal	illegal
illegala	illegal
illinois	illinois
illuminati	illuminati
ilska	anger
image	image
imf	imf
immigranter	immigrants
immunförsvar	immune	immune defense
imperiet	the empire
imperium	empire
import	import
in	in the context: recorded = spela (in)	in
inblandad	mixed
inblandade	involved
inblandning	involvement	incorporation
inbördes	intermutual
inbördeskrig	civil war
inbördeskriget	civil war; civil war	civil war
indelad	divided
indelade	divided	divided into
indelas	divided	categorized
indelat	divided	split
indelning	the subdivision	classification
indelningar	divisions	classifications
indelningen	division	classification
independence	independence
index	index
indian	indian
indiana	indiana
indianer	indians
indianerna	the indians	indians
indianska	red indian	native american
indien	india
indiens	india's	indias
indier	indians
indierna	the indians	indians
indikerar	indicates
indirekt	indirect	indirectly
indisk	indian
indiska	indian
individ	individual
individen	the individual
individens	individual's	the individual's
individer	individuals	subjects
individerna	the individuals
individuella	individual
indoeuropeiska	indo-european
indonesien	indonesia
indonesiska	indonesian
industri	industry	industrial
industrialiserade	industrialized
industrialisering	industrialization
industrialiseringen	indutrialization	industrialization
industriell	industrial
industriella	industrial
industriellt	industrially	industrial
industrier	industries
industrin	industry
infaller	falls
infektion	infection
infektioner	infections	infection
inflation	inflation
inflationen	inflation
influensa	influenza	flue
influensan	the influenza	flu
influensavirus	flu virus	flue virus
influenser	influences
influerad	influenced
influerat	influenced
inflytande	influence
inflytandet	the influence
inflytelserika	influential
information	information
informationen	the information
infrastruktur	infrastructure
infrastrukturen	infrastructure
infödda	native	natives
inför	before
införa	introduce
införande	introduction
införandet	the introduction
införde	introduced
infördes	introduced
infört	introduced
införts	been inserted	introduced
inga	not	no
ingen	no
ingenjör	engineering	engineer
ingenting	nothing
inget	no
ingick	were included
ingmar	ingmar
ingredienser	ingredient	the ingredients	ingredients
ingrid	ingrid
ingripa	interfere	act
ingripande	negative	intervention
ingvar	ingvar
ingå	be a part	be included in
ingående	enter into	in depth
ingår	is
ingått	been part of	entered	entered into
inhemsk	domestic	native
inhemska	native
initiativ	initiative
inkluderade	included
inkluderar	include	includes
inkluderas	is included
inkluderat	included	including
inklusive	including
inkomst	income
inkomster	revenue	income
inkomsterna	the incomes	revenue
inkomstkälla	was added to cold
inlandet	inland	the inland
inleda	initiate
inledande	initial
inledde	started	launched
inleddes	started	began	initiated
inleder	initiates
inledning	introduction	the beginning
inledningen	the beginning	the introduction
inledningsvis	initially	by way of introduction	in the beginning
inleds	starts
inlett	started
inletts	started	initiation
inlägg	post
inlärning	learning
innan	before
innanför	inside	within
inne	inside	in
innebandy	floorball
innebar	was; meant; entailed
inneburit	resulted	meant
innebär	means	mean
innebära	mean
innebörd	meaning
innebörden	meaning	the significance
innefattar	includes
innehade	possessed
innehar	holds
innehas	held	occupied
innehav	owning
innehåll	content
innehålla	include	contain
innehållande	including
innehåller	include	contains
innehållet	content	contents
innehöll	include
innersta	innermost
innerstaden	inner city
inom	within
inre	inner
inrikes	domestic
inriktad	focused on	intent
inriktade	oriented
inriktning	direction	orientation	alignment
inriktningar	direction
inrättades	established	were implemented
insats	contribution	stake
insatser	action
insekter	insects
inser	recognize	realizes
insikt	insight	recognition
inslag	elements	element
inspelad	recorded
inspelning	recording
inspelningar	recordings
inspelningarna	recordings
inspelningen	recording
inspiration	inspiration
inspirerad	inspired
inspirerade	inspired
inspirerades	(was) inspired
inspirerat	inspired
instabil	unstable
installera	install
instiftade	created
institut	institute	institution
institutet	institute
institutioner	institutions
institutionerna	institutions
instruktioner	instructions
instrument	intrument
inställning	attitude	view
insulin	insulin
insåg	realized
inta	taken
intag	intake
inte	not
integration	integration
integritet	integrity
intellektuella	intellectuals	intellectual
intensiv	intensity	intense
intensiva	intensive	intense
intensivt	intensive
inter	inter
interaktion	the interaction	interaction
interna	internal
international	international
internationell	international
internationella	international
internationellt	international	internationally
internet	internet
interstellära	interstellar
intervju	interview
intervjuer	interviews
intet	nothing	no
intill	beside	adjacent to
intog	occupied	seized
intogs	was taken	was captured
intressant	interestingly
intressanta	interesting
intresse	interest
intressen	interests
intresserad	interested
intresserade	interested
intresset	interests	the interest	interest
introducerade	introduced
introducerades	introduced
intryck	impression
inträde	entry
inträffade	occurred	happened
inträffar	occur
intäkter	incomes
intäkterna	the revenues	the revenue
intåg	entry	advent
inuti	inside
invadera	invade
invaderade	invaded
invaldes	was elected
invandrade	immigrated	immigrant
invandrare	immigrants	immigrant
invandring	immigration
invasion	invasion
invasionen	the invasion
inverkan	impact	influence	effect
investeringar	investments
invigdes	inaugurated
invigningen	inauguration	the opening
invånare	resident (-s)	inhabitants
invånarna	inhabitatants; citizens'
inåt	inwards	inwardly
ip	ip
irak	iraq
irakiska	iraqi	irakish
irakkriget	iraq war
iraks	iraq
iran	iran
irans	iran's
iranska	iranian
irland	irland	ireland
irländska	irish
isberg	ice berg	iceberg
isbn	isbn
isen	the ice
ishockey	ice hockey
ishockeyspelare	ice hockey player	hockey players
islam	islam
islamisk	islamic
islamiska	islamic
islamistiska	islamic	islamist
islams	islams	islam's
island	icelandic
isländska	icelandic
iso	iso
isolerad	isolation	isolated
isolerade	isolated
isolering	isolation
isotoper	isotopes
israel	israel	israeli
israelisk	israeli
israeliska	israeli	isrealic
israels	israels	israel's
istanbul	istanbul
istiden	ice age	the ice age
istället	instead
isär	ice	apart
italien	italy
italiens	italy's
italiensk	italian
italienska	italian
iu	iu
ivan	ivan
ivar	ivar
iväg	away
ix	4	the ninth
ja	yes
jack	jack
jackie	jackie
jackson	jackson
jacksons	jackson's	jacksons
jacob	jacob
jacques	jacques
jag	i
jaga	course	hunt	chase
jagar	hunting
jah	jah
jakob	jakob
jakt	hunt	hunting
jakten	the hunt	hunt
jamaica	jamaica
jamaicanska	jamaican
jamaicas	jamaicas	jamaica's
james	james
jan	jan	january
janeiro	janeiro
januari	january
janukovytj	janukovytj
japan	japan
japanerna	japanese
japans	japans	japan's
japansk	japansk	japanese
japanska	japanese
jarl	earl	jarl
jason	jason
java	java
jazz	jazz
jean	jean
jeff	jeff
jefferson	jefferson
jehovas	jehovas	jehova's
jennifer	jennifer
jenny	jenny
jens	jens
jensen	jensen
jersey	jersey
jerusalem	jerusalem
jerusalems	jerusalem's
jesu	jesu
jesus	jesus
jihad	johad	jihad
jim	jim
jimi	jimi
jimmy	jimmy
joachim	joachim
joakim	joakim
joan	joan
jobb	job
jobba	work
jobbade	worked
jobbar	work
jobbet	work	the job
joe	joe
joel	joel
joey	joey
johann	johann	john
johannes	johannes
johans	johan's	johan
johansson	johansson
johanssons	johanssons
john	john
johnny	johny	johnny
johnson	johnson
joker	joker
jolie	jolie	jolies
jon	jon
jonas	jonas
jonatan	jonatan	jonathan
jonathan	jonathan
jones	jones
jonsson	jonsson
jord	earth
jordanien	jordan
jordbruk	agricultural
jordbruket	agriculture	the agriculture
jordbävning	earthquake
jordbävningar	earthquakes
jordbävningen	the earthquake
jorden	the earth	earth	earth; earth; underground
jordens	earth
jorderosion	earth erosion	soil erosion
jordskorpan	earth's crust	earth crust	the earth's crust
jordytan	earth's surface	earth crust
jorge	jorge
josef	josef
joseph	joseph
josé	jose
journal	journal
journalist	journalist
journalisten	the journalist
journalister	journalists
jr	junior
ju	the
juan	juan
judar	jews
judarna	jews
judarnas	jews
judas	judas
jude	jew
judendom	judaism	jewism
judendomen	the judaism	judaism
judisk	jewish
judiska	jewish
judy	judy
jugoslavien	yugoslavia
jugoslaviska	jugoslavian	yugoslavian
jul	christmas
julafton	chistmas eve	christmas eve
juldagen	christmas day
julen	christmas
jules	jules
juli	july
julia	julia
julian	julian
julie	julie
julius	julius
juni	june
junior	junior
jupiter	jupiter
jupiters	jupiter's
juridik	law
juridisk	legal
juridiska	juridical	legal
juridiskt	legally	juridical	judicial
juryn	the jury
juryns	the jury's
jussi	jussi
just	currently	just
justice	justice
juventus	juventus
jämför	compare
jämföra	compare
jämföras	compared
jämförelse	comparison
jämförelser	comparison
jämförelsevis	in comparison	comparatively
jämfört	compared to last	compared	compared (to)
jämlikhet	equality
jämna	even
jämnt	even	evenly
jämte	next (to)	plus
järn	iron	kon
järnmalm	iron ore
järnväg	railroad	rail	railway
järnvägar	failways	railways
järnvägarna	the railways	railways
järnvägen	railroad
järnvägsnätet	railroad network	rail
jönköping	jönköping	jonkoping
jönköpings	jönköpings
jönsson	jönsson	johnsson
jönssonligan	jönssonligan	jonssonligan
kaffe	coffee
kaffet	the coffee
kairo	cairo
kalender	calendar	calender
kalendern	calender
kalifornien	california
kalksten	limestone
kall	cold
kalla	cold
kallad	know as	called
kallade	called
kallades	was called	summoned
kallar	calls
kallare	colder
kallas	called
kallat	called
kallats	was called	called
kallblod	cold blood	cold blooded	draught horse
kalle	kalle
kallt	cold	coldly
kalmar	kalmar
kammare	chamber
kammaren	chamber	the chamber
kamp	struggle	fight
kampanil	kampanil	bell tower	bellfry; bell tower	campanile
kampanj	campaign
kampanjen	campaign
kampen	the struggle	the fight	fight
kampf	kampf
kamprad	kamprad
kan	can be
kanada	canada
kanadas	canada's
kanadensiska	canadian
kanal	channel
kanalen	the channel	channel
kanaler	channels
kanarieöarna	canary islands	the canary islands
kandidat	candidate
kandidater	candidates
kanske	may
kant	kant	edge
kantoner	cantons
kantonerna	the cantons	cantons
kaos	chaos
kap	chapter	cape
kapacitet	the capacity	capacity
kapital	capital
kapitalet	the capital
kapitalism	capitalism
kapitalismen	capitalism
kapitalismens	capitalism's	capitalism
kapitalistiska	capitalistic	capitalist
kapitel	chapter
kapitulation	surrender	capitulation
kapitulerade	surrendered
kapten	captain
karakteristiska	characteristic
karaktär	character
karaktären	the character	character
karaktärer	characters
karaktäriseras	characterizes	is characterised
kardinal	cardinal
karibiska	caribbean
karin	karin
karl	karl
karlsson	karlsson
karlstad	karlstad	phoenix
karlstads	karlstad's
karma	karma
karolinska	karolinska (institute for medicine)	caroline
karriär	career
karriären	career	the career
karta	map	maps
kartan	the map
kartor	maps
kaspiska	caspian
kasta	throw
kastar	throws
katalanska	catalan
katalonien	catalonia
katastrofen	catastrophy	the catastrophy
katastrofer	catastrophes	disasters
kate	kate
kategori	category
kategoriasiens	category of asia
kategoribrittiska	category: british
kategorier	categories
kategorieuropas	category europe
kategorifiktiva	category fictitious
kategorifödda	category: born
kategorikrigsåret	category war years
kategorikvinnor	category women
kategoriledamöter	category: members
kategorimusik	category music
kategorimän	category: men
kategorin	category	the category
kategoriorter	category visited
kategoripersoner	category of persons
kategorirock	category:rock
kategorispelare	category player
kategorisvenska	category: swedish
kategorisvenskar	category swedes
kategorityska	category: german
katekes	catechism
katla	katla (fictive dragon in the classic "bröderna lejonhjärta")
katolicismen	catholisism	catholicism
katoliker	catholics
katolsk	catholic
katolska	catholic
katt	cat
kattdjur	cat	felidae
katten	the cat
katter	cats
kazakstan	kazakstan	kazakhstan
kedja	chain
kedjan	the chain
kedjor	chains
keith	keith
kejsar	emperor
kejsardömet	empire
kejsare	emperor
kejsaren	the emperor
kejsarens	the emperor's	emperors
kejserliga	imperially	imperial
keltiska	celtic
kemi	chemistry
kemikalier	chemicals
kemisk	chemical
kemiska	chemical
kemiskt	chemically
ken	ken
kennedy	kennedy
kenneth	kenneth
kenny	kenny
kent	kent
kenya	kenya
keramik	ceramic	ceramics
kevin	kevin
kids	kids
kiev	kiev
kill	kill
kille	guy
kilometer	kilometer	kilometers
kim	kim
kina	china
kinas	chinas
kinesisk	chinese
kinesiska	chinese
kings	king's
kingston	kingston
kirsten	kirsten	kristen
kiss	kiss
kjell	kjell
kl	hr	at
klan	clan
klar	done
klara	clear
klarade	passed
klarar	do	handle
klart	finished	done
klass	grade; class
klassas	classified
klassen	the class
klasser	classes
klassificera	classifying	classify
klassificeras	classified
klassificering	classification
klassiker	classic
klassisk	classic
klassiska	classic
klassiskt	classical	classic
klaviatur	keyboard
klimat	climate
klimatet	environment	climate
klimatologi	klimatology	climatology	climateology
klippa	cut
klippiga	rocky
klitoris	clitoris
klockan	clock	o'clock
klorofyll	cholophyll
kloster	monastery
klp	klp
klubb	club
klubbar	clubs
klubbarna	clubs	the clubs
klubben	club
klubbens	club
klubblag	club teams
klädd	clothed	coated
kläder	clothes
klädsel	cover
km	kilometers
km²	square kilometre	km2
knapp	scarce	bare
knappast	hardly
knappt	barely
knight	knight
knut	knut	knot
knuten	tied to	bound
knutna	associated	tied
knutpunkt	hub
knutsson	knutsson
knyta	tie
knä	knees	knee
knäppupp	knäppup	knäppupp
ko	co	cow
koalition	coalition
koden	the code
koenigsegg	koenigsegg
koffein	caffein
kognitiv	cognitive
kognitiva	cognitive
kokain	cocaine	cocain
kokpunkt	boiling point
kol	coal; charcoal
koldioxid	co
kolhydrater	carbons	carbohydrates
kollaps	collapse
kollapsade	collapsed
kollektiv	collective	public
kollektivtrafik	public transport
koloni	colony
koloniala	colonial
kolonialism	colonialism
kolonialismen	the colonialism	colonialism
kolonialtiden	the colonial times
kolonier	colonies
kolonierna	colonies
kolonin	colony
koloniserades	is colonized	colonized
koloniseringen	the colonization
kolväten	hydrocarbons	the hydrocarbon
kom	came
koma	coma
kombattant	combatant	combatant; fighter
kombination	combination
kombinationen	the combination	combination
kombinationer	combinations
kombinerad	combined
kombinerade	combined
kombineras	combined
kombinerat	combined
kometer	comets
komiker	comic	comedian
komintern	komintern	comintern
komma	access	get
kommande	upcoming
kommendör	commandor	commander
kommentar	comment
kommentarer	comments
kommenterade	comment	commented
kommer	is
kommersiell	commercial
kommersiella	commercial
kommersiellt	commercial
kommissionen	commission	the commission
kommit	to be	come
kommitté	committee
kommittén	the committee	committee
kommun	municipality
kommunal	communal	municipal
kommunala	local	municipal
kommunen	municipality
kommuner	municipalities	counties
kommunerna	kommunera	municipalities	the municipalities
kommunicera	communicate
kommunicerar	communicates
kommunikation	communications	communication
kommunikationer	communications
kommunism	communism
kommunismen	communism
kommunismens	communism	the communisms	the communism's
kommunister	communists
kommunisterna	communists	communist	the communists
kommunistisk	communistic	communist
kommunistiska	communistic	communist
kommunistpartiet	the communist party
kommunistpartiets	communist party	the communist party	the communist partys
komplett	complete
komplex	komplex	complex
komplexa	complex
komplext	complex
komplicerad	complex	complicated
komplicerat	complicated
komplikationer	complications
komponenter	components
kompositör	composer
kompositörer	composers	compositors
kon	group
koncentration	concentration
koncentrationsläger	concentration camp	concentration camps; kz-camps
koncentrerad	concentrated	concentration
koncentrerade	concentrated
koncept	concept
konflikt	conflict	conflict; strife
konflikten	the conflict	conflict
konflikter	conflicts	conflict
kong	(hong) kong	kong
kongo	congo
kongokinshasa	kong kinshasa	democratic republic of the congo
kongress	congress
kongressen	congress
kongresspartiet	congress party	indian national congress
konkret	concrete
konkreta	concrete
konkurrens	competition
konkurrensen	the competition
konkurrerande	competing
konkurs	bankruptcy
konsekvens	consequence
konsekvenser	consequences
konsekvenserna	consequensis
konsekvent	consistent	consistency
konsensus	consensus
konsert	concert
konserten	the concert	concert
konserter	conserts	concerts
konserterna	the concerts
konserthus	concert hall	concert
konservatism	conservatism
konservatismen	conservatism
konservativ	conservative
konservativa	conservative
konsolen	bracket
konspirationsteorier	conspiracy theories
konst	art
konstant	constant
konstantin	konstantin	constantine
konstantinopel	constantinople
konstaterade	concluded	established	stated
konsten	art	the art
konstitution	constitution
konstitutionell	constitutional
konstitutionella	constitutional
konstitutionen	constitution
konstnär	artist
konstnären	the artist	artist
konstnärer	artists
konstnärlig	artistic
konstnärliga	artistic
konstruerade	constructed
konstruktion	construction
konstverk	work of art	artwork
konsubstantiation	no idea what it means	consubstantion	konsubstantiation	con-substantiation	consubstantiation
konsul	consul	consulting
konsumtion	consumption
konsumtionen	the consumtion	consumption
kontakt	plug	contact
kontaktade	contacted
kontakten	conntact	the contact
kontakter	contact	contacts
kontinent	continent
kontinentala	continental
kontinenten	the continent
kontinentens	the continents
kontinenter	continents
kontinuerlig	continuous
kontinuerligt	continuous	continous
konto	account	sign
kontor	office
kontrakt	agreement	contract
kontraktet	the contract
kontrast	contrast
kontroll	control
kontrollen	control	the control
kontrollera	control
kontrollerade	controlled
kontrollerar	controlling	controls; controlling
kontrolleras	is controlled
kontroverser	controversies
kontroversiell	controversial
kontroversiella	controversial
kontroversiellt	controversial
konung	king
konungarike	kingdom
konungariket	kingdom
konventionella	conventional
konventionen	convention
konventioner	conventions
konvertera	convert	conversion
konverterade	converted
kopia	copy
koppar	copper
koppla	coupling	connect
kopplad	connected to	connected
kopplade	connected
kopplas	connected
kopplat	coupled; connected	connected
koppling	connection
kopplingar	connections
kopplingen	the connection	coupling
koprolali	coprolalia	coporolalia
koranen	the koran	the quran
korea	korea
koreakriget	the korean war
koreanska	korean
korn	korn	barley
korrekt	correct
korrekta	correct
korruption	corruption
korruptionsindex	corruption index
kors	cross
korset	cross
kort	short
korta	short
kortare	shorter
kosmiska	the cosmic	cosmic
kosovo	kosovo
kosovos	kosovo's
kostade	cost
kostar	costs
kostnaden	cost
kostnader	costs	expenses
kostnaderna	costs	the costs
kostym	costume
kr	kronas
kraft	force	power
kraften	the force	power
krafter	forces
kraftfull	forceful	powerful
kraftig	strong
kraftiga	strong	powerful
kraftigare	greater	more powerfully
kraftigt	heavily
kraftverk	power plant
krav	requirement	demands
kraven	the demands	requirements
kravet	requirement	the demand
kreativitet	creativity
krets	sphere	circuit
kretsar	circles
kretsen	the order
krig	war
krigare	warriors	warrior
krigen	the wars	wars
kriget	the war
krigets	the war's
krigsmakt	military power	armed forces
krigsmakten	armed forces
krigsslutet	end of war; war's end	end of the war
kriminella	criminal
kring	around
kris	crisis
krisen	the crisis
kriser	crises
kristen	christian
kristendom	christianity
kristendomen	chritianity	christianity
kristendomens	the christianity's	christianity's
kristi	christ
kristian	kristian
kristiansson	kristiansen
kristinas	kristina's
kristna	christian
kristus	christ
krita	chalk
kriterier	criteria
kriterierna	criteria
kritik	criticism	critisism	critique; criticism
kritiken	criticism	the criticism	the critique
kritiker	critics	critiques
kritikerna	critics	the critics	critiques
kritiserade	critisized	criticized
kritiserades	critisized	critizised
kritiserar	criticize
kritiserat	criticized	criticised
kritiserats	criticized	critized
kritisk	critical
kritiska	critical
kritiskt	critical
kroatien	croatia
kroatiens	croatia's	croatias	croatian
kroatiska	croatian
kromosom	chromosome
kromosomer	chromosomes
kromosomerna	chromosomes	the chromosomes
krona	crown
kronan	crown	kronan
kronisk	chronic
kroniska	chronic
kronor	kronor	crowns
kronprins	crown prince
kronprinsen	crown prince	the crown prince
kronprinsessan	crown princess
kropp	body
kroppar	cells	bodies
kroppen	body	the body
kroppens	the body's	the bodies
krossa	crush
kryddor	spices
kräva	demand
krävde	demanded
krävdes	were required
kräver	requires
krävs	needs
krävt	taken	required
krönika	chronicle
kröntes	crowned
kub	cube
kuba	cuba
kubanska	cuban
kubas	cuba	cuba's
kuben	the cube
kuiperbältet	the kuiper belt	the cuyper belt
kulmen	the acme	peak
kulminerade	culminated
kultur	culture
kulturarv	culture heritage	cultureheritage	cultural heritage
kulturell	cultural
kulturella	cultural
kulturellt	cultural	culturally
kulturen	culture	the culture
kulturer	cultures
kunde	could
kunder	customer
kung	king
kungafamiljen	the royal family
kungahuset	royal family	royal house
kungamakten	monarchy	the monarchy
kungar	kings
kungariket	kingdom	the kingdom
kungarna	the kings
kungen	king	the king
kungens	the king's
kunglig	royal
kungliga	royal
kunna	to	be able
kunnat	could	could have been
kunskap	knowledge
kunskapen	the knowledge	knowledge
kunskaper	knowledge
kupol	cupola	combatant	dome	cu
kupp	kupp	coup (d'etat)
kurder	kurds
kurderna	kurdish
kurdisk	kurdish
kurdiska	kurdish
kurdistan	kurdistan
kurfursten	elector
kuriosa	bric-a-brac	trivia
kurs	course
kurt	kurt
kusin	cousin
kust	coastal	coast
kusten	the coast
kuster	coasts
kusterna	the coasts	coasts
kustlinje	coastline
kuwait	kuwait
kvadratkilometer	square kilometer	square kilometers
kvalificerade	qualifying
kvalitet	quality
kvar	left
kvarstod	remained
kvarstår	remains
kvarter	quarter	block
kvarteret	quarter	the neighborhood
kvartsfinalen	quarter finals	quarterfinals
kvarvarande	remaining	lasting
kvast	broom	groom
kvicksilver	mercury	quicksilver	witty zeal
kvinna	woman
kvinnan	woman
kvinnans	female
kvinnlig	female
kvinnliga	female
kvinnor	female	women
kvinnorna	the women	women
kvinnornas	womens	the women's
kvinnors	women	women's
kväll	evening
kvällen	the evening
kväve	nitrogen
kyla	cold
kyrilliska	cyrillic
kyrka	church
kyrkan	the church
kyrkans	the church's	the churche's
kyrkliga	religious	from the church
kyrkor	churches
kyrkorna	churches	the churches
kyros	cyrus
källa	source
källan	source	kallan	the source
källkod	source code
källor	source
källorna	the sources
kämpa	fight
känd	known	famous
kända	known
kände	felt
känna	known	know
kännedom	knowledge
känner	know
kännetecken	distinction	sign
kännetecknas	is characterized	characterized (by)	characterized
känns	feels
känsla	feeling
känslan	feeling	the feeling
känslig	susceptible
känsliga	1st&2nd: fragile 3rd: sensitive	bilge accordance
känslor	feelings
känt	known	famous
kär	in love
kärlek	love
kärleken	the love
kärna	core
kärnan	core	the core
kärnkraft	nuclear power
kärnkraftverk	nuclear power plant	nuclear powerplant
kärnor	cores	core
kärnvapen	nuclear weapons
köket	cuisine	the kitchen
köln	köln
kön	gender	sex
könen	the sexes	equality
könsorgan	genitals	sex organ
könsorganen	sex organs	the reproductive organs	the genitals
köp	purchase
köpa	purchase	buy
köpenhamn	copenhagen
köpenhamns	copenhagen's
köper	making
köpmän	traders	merchants
köpt	purchased	bought
köpte	purchased	bought
kör	run
köra	run	drive
körberg	körberg
körs	driven	being driven
kött	cones	meat
l	l
la	la
laboratorium	laboratory
ladda	load
laddade	charged
laddning	charge
lade	laid	seized
lades	put	was
ladin	ladin
lag	law
lagar	laws
lagarna	the laws
lagen	the law	law
lager	layer
lagerkvist	lagerkvist
lagerlöf	lagerlof	lagerlöf
laget	the team	stroke
lagets	the team's	substrate
lagförslag	bill	lagforslag
lagliga	legal
lagras	stored
lagring	storage
lagstiftande	legislative	legislating	legislation
lagstiftning	law-making
lagstiftningen	law-making	legislation
lagt	laid	added
lagts	added
laila	laila
lake	lake
land	country
landet	the country
landets	the country's	its
landområden	land areas	land
lands	on land
landsbygden	rural area
landshövding	county governor	governor
landskap	province	landscape
landskapen	the landscapes	landscapes	landscape
landskapet	landscape
landskommun	rural municipality
landslag	national team
landslaget	the national team
landsting	county	county council
lanka	lanka	(sri) lanka
lanserade	introduced	launched
lanserades	launched	was launched
lanseringen	the release	launch
laos	laos
larry	larry
lars	lars
larsson	larsson
larssons	larsson's
laryngoskop	laryngoscopes	laryngoscopy	llaryngoscope	laryngoscope
lasse	lasse
lastbilar	truck	trucks
lat	methacrylate
latin	latin
latinamerika	latin america
latinamerikanska	latin-american	latin american
latinet	latin
latinets	the latin	the latin's
latinska	latin
laura	laura
lava	lava
lawrence	lawrence
le	smile
led	suffered
leda	lead
ledamot	member	representative
ledamöter	commissioners
ledamöterna	the commissioners	commisioners	the members
ledande	conductive	leading
ledare	conductors	leader
ledaren	leader
ledarna	the leaders	conductors
ledarskap	leadership
ledda	run (by)
ledde	led
leddes	passed	was led
leden	hinge	lines	the route
leder	leads	leading (to)	lead
ledger	ledger
ledning	guidance
ledningen	the lead
leds	led by	passed
lee	lee
leeds	leeds
left|px	left px
legat	layed
legend	legend
legenden	legend
legender	legends
legitimitet	legitimacy
leipzig	leipzig	liepzig
lejon	lion
lejonet	the lion
lena	lena
lenin	lenin
lenins	lenin's
lennart	lennart
lennon	lennon
leo	leo
leonard	leonard
leonardo	leonardo
leopold	leopold
les	les
let	cleanly
leta	search
lett	led (to)
lettland	latvia
leukemi	leukemia
lev	lev
leva	live
levande	live
levde	lived
lever	living	live
levern	the liver
levnadsstandard	living standard	standard of living
levnadsstandarden	the standard of living	living standard
levt	survived
lewis	lewis
lexikon	lexicon
liam	liam
libanon	lebanon
liberala	liberal
liberaler	liberals
liberalism	liberalism
liberalismen	the liberalism
liberty	liberty
library	library
libyen	libya
lida	sheath	suffer
lidande	sufferer
lider	suffers
lidit	suffered
liechtenstein	liechtenstein
life	life
liga	league
ligacupen	league cup
ligan	league
ligga	lies, lie	lie
liggande	lie	placed
ligger	lies
light	light
lik	similar	alike
lika	similar	equal	alike
likartade	similiar	similar
likaså	also	as well
likhet	similar	resemblance	like
likheter	similarities	similarity
liknade	similar	looked like
liknande	similiar	similar
liknar	similar
liknas	compared to	likened
liksom	and	as is
likt	like
likväl	nevertheless	still	as well
likör	cordial	liqueur	liqeur	liquor	liquer
lilla	small
lima	lima
lina	line	lina
lincoln	lincoln
linda	linda
lindgren	lindgren
lindgrens	lindgren's	lindgren	lindgrens
lindh	lindh
linje	line
linjen	the line
linjer	routes	lines
linjerna	the lines	lines
linköping	linköping
linköpings	linkopingas	linköping's
linné	linneus
linux	linux
lisa	lisa
lisbet	lisbet
lissabon	lisbon
lissabonfördraget	treaty of lisbon	lisbon treaty
list	cunning
lista	list
listade	listed
listan	the list
listor	lists
listorna	menus	the lists
litauen	lithuania
lite	little
liten	small
liter	liters
litet	small
litteratur	litterature
litteraturen	literature
litterär	literary
litterära	literary	literal
liv	life
livealbum	live album
liverpool	liverpool
liverpools	liverpool's
livet	the life	life
livets	life's	the life's
livslängd	life	life expectancy
livsmedel	food
livsstil	life style	lifestyle
livstid	lifetime
liza	liza
ljud	sounds	noise
ljudet	the sound	noise
ljung	heather
ljungström	ljungström
ljus	light
ljusare	brighter	lighter
ljuset	the light	light
locka	tempt
lockar	attracts	curls
locke	locke
loggbok	journal	log book	logbook	log
logik	logic
logotyp	logotype
lois	lois
lojalitet	loyality
lokal	local
lokala	local
lokaler	studios	place
lokalt	locally	local
london	london
londons	london's
lopp	course, passage	race
loppet	the race
lord	lord
loss	unstuck	off
lost	lost
lotta	lotta
louis	louis
louise	louise
louisiana	louisiana
lovade	promised
lovat	promised
lp	lp
lsd	lsd
lucas	lucas
lucia	lucia
lucky	lucky
ludvig	louis	ludvig
ludwig	lugwig	ludwig
luft	air
luften	air
lugn	calm
lugna	calm
lukas	lukas
luleå	luleå
luminositet	luminosity
lundell	lundell
lundgren	lundgren
lunds	lund's
lunginflammation	pneumonia
lungorna	the lungs
lupus	lupus
lust	desire
luther	luther
luthers	luthers	luther's	luther
lutherska	lutheran
lutning	closing	angle	incline
luxemburg	luxemburg
lycka	happiness
lyckade	successful
lyckades	succeeded
lyckan	the happiness	happiness
lyckas	succeed
lyckats	succeeded
lyder	reads	obeys
lyfta	lift
lyfter	lift	lifts	lifting
lyrik	poetry
lysande	brilliant
lyssna	listening	listen
lyssnade	listened
lyssnar	listens	listen
läge	location	mode
lägenhet	apartment	appartment
läger	camp
läget	position	location
lägga	put	lay
läggas	laid
lägger	put	lies
läggs	put before; submitted; put	lay
lägre	lower
lägret	the camp	camp
lägst	lowest	lowermost
lägsta	lowest
läkare	doctor	doctors
läkaren	the doctor
läkemedel	medicine	drugs
läkemedelsverket	medicines work	medical products agency
lämna	leave
lämnade	left
lämnades	left
lämnar	leaves
lämnas	left
lämnat	left
lämningar	remains	remnants
lämplig	suitable
lämpliga	suitable
lämpligt	suitable
län	state
länder	states	countries
länderna	the countries
ländernas	the countries	countries
länders	countries'	countrie's
längd	length
längden	the length	length	lenght
länge	long
längre	longer
längs	along
längst	longest	farthest
längsta	longest	maximum
längtan	longing
länk	link
länkar	links
läns	county	county's
lär	teach	learn
lära	lara	learn	get to know
läran	teaching	the teaching
lärare	teacher
lärda	literate	savants
lärde	learned
lärjungar	disciples	disciple
läror	teachings
lärt	learned	learnt
läs	read
läsa	read
läsare	reader	readers
läsaren	the reader
läser	read	are reading
läses	read	is read
läsning	reading
läst	read	load
läste	read
lät	made	had
lätt	easy
lätta	light	lighten
lättare	easier
låg	low
låga	low
lågt	low
lån	loan
låna	borrow	lana
lånat	borrowed
lång	long
långa	long
långbåge	longbow	long arc	long bow	langbage
långfilm	feature film	feature movie
långhårig	rough	long haired	long-haired
långsamma	slow
långsammare	slower
långsamt	slowly
långt	far
långtgående	far-reaching
långvarig	of long duration	prolonged; lengthy; long	long
långvariga	long-standing
långvarigt	long-running	prolonged	long-standing
låt	song
låta	let
låtar	songs
låtarna	the songs
låten	the song
låter	let
låtit	let	ordered
låtskrivare	song writers
löfte	promise
löften	promises
lön	salary	wage; salary
löner	salaries
lönneberga	lönneberga	lonneberga
löpande	running	assembly	conveyor (belt)
löper	runs
lördagen	the saturday	saturday
lösa	solve
lösas	solved
löser	solves
lösning	solution	solution; resolution
lösningar	solutions
lösningen	the solution	solution
lösningsmedel	solvent
löst	solved	1st sentence: loosely; 2nd & 3rd: solved
löstes	solved
mabel	mabel
machu	machu
madagaskar	madagascar
madeira	madeira
madeleine	madeleine
madonna	madonna
madrid	madrid
maffia	mob	mafia	the mob
maffian	mafia
magdalena	magdalena
magic	magic
magnetfält	magnetic	magnetic field
magnetiska	magnetic
magnitud	magnitude
magnus	magnus
magnusson	magnusson
mahatma	mahatma
maiden	maiden
maidens	maidens
main	main
maj	may
majoritet	majority
majoriteten	the majority
majs	corn
makadam	tarmac	metal	macadam
make	husband
makedonien	macedonia
makedonska	macedonian	makedonish
makt	power
makten	the power
maktens	the powers	the power's
makter	powers
malaysia	malaysia
malcolm	malcolm
malin	malin
malmö	malmö	malmo
malmös	malmö's
malta	malta
mamma	mother
man	one
manager	manager
manchester	manchester
mandat	mandate
mandatperiod	term	term (of office)	term of office
mandelas	mandelas	mandela's
mando	command
manhattan	manhattan
mani	mani	mania
maniska	manic	maniac
mankell	mankell
manlig	male	manly
manliga	male
mannen	art	the man
mannens	man	man's
mans	man's
manson	manson
manteln	the mantle
manuel	manuel
manus	script
manuskript	script
mao	mao
maos	maos	mao's
marco	marco
marcus	marcus
margaret	margaret
maria	maria
marie	marie
mariette	mariette
marijuana	marijuana
marilyn	marilyn
marina	marina	marine
marinen	navy	marines
marino	marino
mario	mario
marissa	marissa
mark	ground, soil, territory	ground
markant	considerably	marked
marken	soil
markera	mark
markerade	selected	marked
markerar	selects	marks
marklund	marklund
marknad	market
marknaden	the market	market
marknader	markets
marknadsekonomi	market economy
markus	marcus
marley	marley
marleys	marley's
marocko	morocco	marocco
mars	march
marshall	marshall
martin	martin
marx	marx
marxism	marxism
marxismen	marxism	the marxism
marxistisk	marxist	marxistic
marxistiska	marxist
mary	mary
maskiner	machines
massa	mass
massachusetts	massachussetts	massachusetts
massakern	massacre
massan	mass
massiv	massive
massiva	solid	massive
massmedia	media	mass media
massor	lots	(in) masses
master	master
mat	food
match	game	match
matchen	the game	match
matcher	matches	games
matcherna	the games	games
matematik	mathematic	mathematics
matematiken	mathematics
matematiker	mathematician
matematisk	mathematical	mathematic
matematiska	mathematical
maten	the food
materia	matter	materia
material	material
materialet	the material	material
materiella	material
matrix	matrix
mats	mat's
matt	matt
matteus	matthew	matteus
matteusevangeliet	gospel of matthew	book of matthew
matthew	matthew
mattias	mattias
mattis	mattis
maurice	maurice
max	max
maya	maya
med	with
medan	while
medarbetare	employees	coworker
medborgare	citizens
medborgarna	the citizens	citizens
medborgarskap	citizenship
medborgerliga	civil
meddelade	informed; announced	stated
meddelande	message
meddelanden	messages
medel	middle	medium
medelhavet	mediterranean sea
medelhavsklimat	mediterranean climate
medelhavsområdet	the mediterranean region	the mediterranean area
medelklassen	middle class
medellivslängd	average lifespan	life expectancy
medeltemperaturen	median temperature	the average temperature
medeltid	the medieval times
medeltida	middleaged	medival
medeltiden	middle ages
medeltidens	medieval
medelålder	middle age
medför	entails	result
medföra	bring	lead; result in, imply; entail	result
medförde	brought	resulted
medfört	resulted	led to
media	media
medicin	medicine
mediciner	medicines
medicinering	medication
medicinsk	medical
medicinska	medicinal	medical
medicinskt	medical
medier	media	medias
mediet	medium	the medium
medina	medina
medlem	member
medlemmar	members
medlemmarna	members	the members
medlemskap	membership
medlemsstat	member state
medlemsstater	member states	member-state
medlemsstaterna	member	member states
medlemsstaternas	member state	member states
medverka	take part	participate
medverkade	participated; contributed	participated
medverkan	the contribution
medverkar	contribute	contributes
medverkat	participated
medvetande	awareness	consciousness
medveten	conscious	aware
medvetet	consciously
medvetna	aware
mekaniska	mechanical
mekka	mecka
melankoli	melancholy
melker	melker
mellan	between
mellanfot	metatarsals	metatarsus	metatarsal	metatarsal bones
mellankrigstiden	interwar years	interwar period
mellanrum	gap	space
mellanöstern	the middle east	middle east
mellersta	middle	the middle
melodier	melodies
melodifestivalen	eurovision song contest
memoarer	memoirs
memorial	memorial
men	but
menade	meant
menar	means
menas	means
menat	meant
mengele	mengele
mening	meanings	sentence
meningar	sentences
mental	mental
mentala	mental	mentala
mer	more
mera	more
mercurys	mercury's	mercurys
merkurius	mercury
merparten	most	the majority	larger part
merry	merry
mesopotamien	mesopotamia
messi	messi
messias	messiah
mest	mostly
mesta	most
mestadels	mostly
metabolism	metabolism
metaforer	metaphores	metaphors
metall	metal
metaller	metals
metallica	metallica
metan	methane
meter	metre	meter
metionin	methione	methionine
metod	method
metoden	the method
metoder	methods
metro	metro
mexico	mexico
mexikanska	mexican
mexiko	mexico
meyer	meyer
mfl	etc	etc.
miami	miami
michael	michael
michail	michail
michel	michel
michelle	michelle
michigan	michigan
mick	mike (microphone)
microsoft	microsoft
midsommar	midsummer
mig	me
miguel	miguel
mikael	mikael
mike	micke	mike
mil	mile	swedish miles	mil
milan	milan
milano	milano
mild	mild
milda	mild
mildare	cooler	milder
miley	miley
militär	military
militära	military
militären	the military
militärer	soldiers
militärt	military	militarily
miljard	billion
miljarder	billions
miljon	million
miljoner	milions	millions
miljontals	millions
miljö	environment
miljöer	environment	environments
miljön	environment	the environment
miljöproblem	environmental problem	environmental problems
miller	miller
milt	mild
min	my
mina	mine
mind	mind
mindre	smaller	less
mineral	mineral
mineraler	minerals
miniatyr	miniature
miniatyr|	miniature
miniatyr|en	thumbnail
miniatyr|karta	thumbnail map	miniature|map
miniatyr|px|den	miniature
miniatyr|px|en	miniature
miniatyr|px|ett	miniature
minister	minister
ministerrådet	minister counsellor
ministrar	ministers
minne	memory
minnen	memories	memory
minnet	the memory	memory
minns	remembers	remember
minoritet	minority
minoriteten	minority
minoriteter	minorities
minoritetsspråk	minority language
minska	reducing	reduce
minskad	decreased	reduced
minskade	was reduced
minskar	decrease	diminishing
minskat	decreased	has decreased	reduced
minskning	decline	decrease
minst	at least
minsta	minimum
minut	minute
minuter	minutes
miss	miss
missbruk	addiction	abuse
missförstånd	misunderstanding
misshandel	assault	abuse
mission	mission
missionärer	missioners	missioner
misslyckade	failed
misslyckades	failed
misslyckande	failure
misslyckas	fail	fails
misslyckats	failed
missnöje	dissatisfaction
missnöjet	grievance	discontent
misstag	mistake
misstänkt	accused	suspect	suspected of
misstänkta	suspected	suspect
mitt	my	center
mitten	middle
mix	mix
mjölk	milk
mm	millimeter	etc.
moberg	moberg
mod	courage	mod
mode	fashion
modell	model
modellen	the model
modeller	models
moder	mother
moderata	moderates	moderate
moderaterna	the moderate	the moderates	moderates
modern	modern
moderna	modern
modernare	mor modern	more modern
modernismen	modernism
modernistiska	modernistic
modernt	modern
modersmål	native language	mother tongue
modet	the fashion	fashion
modo	modo
mohammed	mohammed
moldavien	moldova
molekyler	molecules
moln	cloud
mona	mona
monaco	monaco
monark	monarch
monarken	the monarch	monarch
monarki	monarchy
monarkin	the monarchy
monetära	monetary
mongoliet	mongolia
monica	monica
monicas	monica	monica's
monografi	thesis	monography	monograph
monopol	monopoly
monoteism	monotheism
monoteistiska	monotheistic
monroe	monroe - it's a persons name	monroe
monster	monster
montana	montana
monte	assembly
montenegro	montenergo	montenegro
monument	monument
moore	moore
mor	mother
mora	mora
moral	morality
moralisk	moralic	moral
moraliska	moral
moraliskt	morally
mord	murder
morden	murders	the murders
mordet	the murder
morgan	morgan
morgon	morning
morgonen	the morning	am
morris	morris
moseboken	genesis
moses	moses
moskva	moscow
mot	against
motion	motion
motiv	subjects	motif
motiveringen	the motivation
motivet	the motive
motor	engine
motors	engine's
motorväg	freeway	high way	motorway	highway	interstate
motorvägar	highways
motorvägarna	the highways
motorvägen	motorway	highway
motsats	contrary
motsatsen	the opposite	opposite
motsatt	opposite
motsatta	opposite
motsatte	opposed
motstånd	resistance	opposition
motståndare	opponents
motståndaren	the opponent	adversary
motståndarna	the opponents	opponents
motståndet	the resistance	the resistence
motståndsrörelsen	the resistance
motsvarande	corresponding to	corresponding
motsvarar	comparable	corresponds
motsvarighet	equivalent
motsättningar	oppositions	frictions; clashes
mottagande	host	reception
mottagare	recipient	receiver
mottagaren	the receiver	the recipient
mottagarens	the reciever	the receivers	the receiver's
motto	motto
mottog	received
motverka	prevent	counteract
mountain	mountain
movie	movie
mozart	mozart
mozarts	mozart's
moçambique	mozambique
mr	herr	mr
ms	motor ship
mtv	mtv
muhammad	muhammad
muhammed	muhammed
muhammeds	mohammed's	muhammed's
mullusfiskar	mullets	don't know what it is except for a kind of fish	goatfish	mullusfiskar	red mullet	mullet	goatfishes
mun	oral	mouth
munnen	the mouth	mouth
mur	wall
muren	wall
murray	murray
muse	muse
museer	museums
museet	the museum
museum	museum
music	music
musik	music
musikalen	the musical
musikalisk	musical
musikaliska	musical
musikaliskt	musically talented	musical	musically
musiken	the music
musikens	the music's
musiker	musicians	musicants
musikstil	music still	music style
musikstilar	music genres	music
musikvideo	music video
musikvideon	music video
musikvideor	music videos
muskler	muscles
musklerna	muscles	the muscles
muslim	muslim
muslimer	muslims
muslimerna	muslims	the muslims
muslimsk	muslim; muslem	muslim
muslimska	muslim
mussolini	mussolini	mossolini
mussolinis	mussolini's
mutationer	mutations
mycket	very	much
myndighet	authoroty	authority
myndigheten	the authority
myndigheter	authorities
myndigheterna	authorities	the authorities	the authoroties
mynnar	opening
mynning	outfall	muzzle	mouth
mynt	coins	coin
myntade	coined
myntades	coined	was coined
mysterium	mystery
mystiska	mystical
myter	myths
mytologi	mythology
mytologin	mythology
mytologiska	mytholigical	mythological
mäktiga	powerful
mäktigaste	powerful	most powerful
mälaren	mälaren
män	men
mängd	volume	amount
mängden	amount	the amount
mängder	amounts	amount
männen	the men	men
människa	man
människan	the human	people
människans	humans	mankinds	human
människas	human's; man's	human
människor	human	people
människorna	men	the humans
människors	humans	people's
mänsklig	human
mänskliga	human
mänskligheten	humanity
mänsklighetens	humanity's	humanities
mänskligt	human
märke	badge	label
märken	brands	sign
märks	labeled	notice	noted
märktes	labeled
märta	märta
mästare	master
mästarna	the champions	the masters
mäta	compare	feeding
mäter	measuring	measure
mätningar	measurements	measurments
mäts	measured	is measured
mätt	measured	dull
må	feel	may
mål	case	mal
måla	target
målade	painted
målare	grinders	painter
målen	goals
måleri	painting
målet	the target
målning	painting
målningar	paintings
målningen	milling	the painting
målvakt	goalee	goalkeeper
målvakten	the goalkeeper
mån	concerned
månad	month
månaden	the month	months	month
månader	months
månaderna	months
månar	moons
månarna	moons
måne	moon
månen	the moon	man
månens	the moon's	the moons
många	many
mångfald	diversity	variety
måste	have to	must
mått	measurement	measure
möjlig	possible
möjliga	possible
möjligen	possibly
möjliggjorde	made possible	allowed
möjliggör	enables
möjlighet	oppertunity	possibility
möjligheten	the possibility
möjligheterna	possibilities	the possibilities
möjligt	possible
mönster	marks
mördad	murdered	murderd
mördade	murdered
mördades	murdered	was murdered	murder was
mörk	dark
mörkare	darkey	darker
mörker	dark	darkness
mörkt	dark
möta	meet
möte	meeting
möten	meetings
möter	meets	meet
mötet	the meeting
mötley	mötley
möts	meet	meets
mött	faced	met
mötte	motte	met
möttes	met
münchen	munchen	munich
n	n
nacka	nacka
nagasaki	nagasaki
namibia	namibia
namn	name
namnen	the names	names
namnet	name	the name
nancy	nancy
napoleon	napoleon
napoleons	napoleon's
narkotika	narcotics
nasa	nasa
nash	nash
nathan	nathan
nation	nation
national	national
nationalencyklopedin	the national encyclopedia
nationalförsamlingen	national assembly
nationalism	nationalism
nationalismen	nationalism
nationalister	nationalists
nationalistiska	nationalistic
nationalitet	nationality
nationalpark	national park
nationalparker	national parks
nationell	national
nationella	national
nationellt	nationally
nationen	the nation
nationens	the nation's	nation
nationer	nations
nationerna	the nations	nations
nationernas	the nation's	the nations
nations	nations
nato	nato
natt	night
natten	overnight
nattetid	overnight
natur	nature
natural	natural
naturen	the nature	nature
naturens	nature's
naturgas	natural gas
naturlig	natural
naturliga	natural
naturligt	natural
naturligtvis	course	naturally
naturresurser	natural resources
naturtillgångar	natural resources
naturvetenskapliga	scientific
nazismen	nazism
nazisterna	nazis
nazisternas	the nazi's	nazi
nazistiska	nazi
nazityskland	nazi germany
nazitysklands	nazi germany's	nazi germany
ned	down	bottom
nedan	below
nederbörd	rainfall	precipitation
nederbörden	precipitation	the precipitation
nederlag	defeat
nederländerna	the netherlands	netherlands
nederländska	netherlands	dutch
nedgång	decline	decreases	fall
nedre	lower
nedsatt	impaired	reduced	decreased; diminished
nedåt	downward	down; downwards
need	need
negativ	negative
negativa	negative
negativt	negative
neil	neil
nej	no
nelson	nelson
neo	neo
neologi	neologism	neology	neologi	a new logical
nepal	nepal
neptunus	neptunes	neptune
ner	bottom
nere	down
nervosa	nervosa
nervsystemet	nervous system	the nervous system
neutral	neutral
neutrala	neutral
neutralitet	neutral
neutralt	neutral
neutroner	neutrons	neutron
nevada	nevada
newport	newport
newton	newton
newtons	newton's
nf	nf
nhl	nhl
ni	you
nickel	nickel
nicklas	niclas	nicklas
niclas	niclas
nietzsche	nietzsche
nietzsches	nietzsche's
nigeria	nigeria
nikki	nikki
niklas	niklas
nikola	nikola
nikolaj	nikolaj	nicholas
nils	nils
nilsson	nilsson
nio	nine
nionde	ninth
nirvana	nirvana
nivå	niva	level
nivåer	levels
nivån	level
nixon	nixon
njurarna	the kidneys
nku	nku
nobel	nobel
nobelkommittén	the nobel commitee
nobelpriset	the nobel prize
nobelpristagare	nobel laureate (-s); nobel prize winner (-s)
nobels	nobel's	nobel
nobelstiftelsen	nobel foundation
nog	sufficiently	enough
noga	carefully
noll	zero
nominerad	nominate	nominated
nominerades	was nominated	nominated
nomineringar	nominations
nord	north
nordafrika	north africa
nordamerika	north america
nordamerikanska	north american
norden	scandinavia; (nordic area; region)	the nordic countries
nordens	the scandinavian countries'	nordic
nordirland	north ireland
nordisk	norse	nordic
nordiska	nordic
nordiskt	nordic
nordkorea	north korea	north koreans
nordkoreanska	north korean
nordkoreas	north coreas
nordliga	northernly	northern
nordligaste	northern	northernmost
nordost	north east	the northeast
nordsjön	north sea
nordväst	north west	northwest
nordvästra	northwest	north western
nordöst	northeast
nordöstra	nordeastern	northeast
norge	norway
norges	norway's
normal	normal
normala	normal
normalt	normally	normal
norman	norman
normer	norms	standards
norr	north
norra	northern
norrköping	norrköping
norrköpings	norrköpings
norrland	northern	norrland
norrlands	northern sweden's	lapland's	norrland
norrmän	norwegians
norrut	north
norsk	norwegian
norska	norwegian
norstedt	norstedt
norstedts	collins	norstedt's
north	north
notation	notation
noter	notes	notation
notera	note
noterade	noted
nou	nou
nova	nova
november	november
now	now
nr	no.	number	no
nsdap	nsdap
nu	now
nuförtiden	nowadays	today
nukleotider	nucleotides	nucleotide
numera	now	nowadays
nummer	number
nutid	present
nutida	present(-day); contemporary
nuvarande	current
ny	new
nya	new
nyare	newer
nybildade	newly formed
nye	new
nyfödda	newborn
nyheten	news
nyheter	news
nyligen	recently
nytt	new
nytta	good	useful
nyval	re-election	new election	election
nämligen	namely
nämnas	mentioned	include
nämnda	said
nämnde	mentioned
nämner	mentions
nämns	mentioned
nämnts	mentioned
när	when
nära	close	near
närhet	closeness
näring	nutrition
näringsliv	business
näringslivet	economic life	industrial life	business
närliggande	adjacent	nearby
närma	approach
närmade	approached
närmar	close in	closing
närmare	close to
närmast	mediately	closest	nearest
närmaste	closest
närstående	relative	relatives	kindred
närvarande	present (-ly)	present
närvaro	attendance
näsan	the nose
näst	second (to)
nästa	next
nästan	almost
nät	web	net(work)
nätet	net	the internet
nätverk	network
nätvingar	natvinger	lacewings	net-winged insects	neuropteran	net wings, it's a animal	neuropterans	neuroptera	nätvingar	netwings	lacewing	natvingar
nå	reach
nåd	mercy	grace
nådde	reached
nåddes	reached
någon	someone	anybody
någonsin	ever
någonstans	somewhere
någonting	anything
någorlunda	fairly	somewhat
något	any	something
några	few	a few
når	reach
nås	reached
nått	reached
nöd	distress
nödvändig	necessary
nödvändiga	necessary	essential
nödvändigt	neccessary	necessary
nödvändigtvis	by necessity	necessarily
nöjd	content
o	oh
oavgjort	draw
oavsett	regardless; whether; irrespective of	regardless
obama	obama
obamas	obama's
obelix	obelix
oberoende	independent
objekt	object
objekten	items	the objects
objektet	the object	object
obligatorisk	obligatory	mandatory
obligatoriskt	mandatory
observationer	observations
observatörer	observers
observera	observe
observeras	observed	is noticed	is observed
oc	oc
oceanen	the ocean
och	and
ocheller	and/or
också	also
ockupation	occupation
ockupationen	the occupation	occupation
ockuperade	occupied
ockuperades	occupied
ockuperat	occupied
oden	oden
odens	odin's	oden's
odlade	grew
odlas	cultured
odling	cultivation
oecd	oecd
oerhörd	tremendous
oerhört	tremendously
of	av
off	off
offensiven	offensive	the offensive
offentlig	public
offentliga	public
offentligt	public	publicly
offer	victim
office	office
officerare	officers	officer
official	official
officiell	official	authentic
officiella	official
officiellt	official	officially
offren	victims
offret	the victim	offering
offside	offside
ofta	often
oftare	more often	more
oftast	usually	most often
oförmåga	inability	failure
ogillade	disliked
oklart	clear
oktober	october
oktoberrevolutionen	the october revolution	october revolution
okänd	unknown
okända	unknown
okänt	unknown
ola	ola
olagligt	illegal
olika	different	variety
oliver	olives
olja	oil
olle	olle
ollonet	penis head	glans	the glans
olof	olof
olsson	olsson
olycka	incident	accident	disaster
olyckan	the accident
olyckor	accidents
olympia	olympia
olympiastadion	olympa stadium	olympic stadium
olympiska	olympic
om	of	for	if
ombord	onboard
omedelbar	immediate
omedelbart	immediately	immediate
omfatta	cover
omfattade	included
omfattande	large	massive; extensive
omfattar	encompass
omfattas	comprise	subject
omfattning	extent
omger	surrounds	surrounding the
omges	surrounded
omgivande	surrounding	surounding
omgiven	surrounded
omgivning	surrounding	surroundings	ambient
omgivningen	surroundings	the surrounding	ambient
omgående	immediate
omgångar	in turns; periods; mandates
omgången	round
omkom	perished	died; was killed	died
omkring	surrounding
omkringliggande	surrounding	neighbouring
omloppsbana	orbit
omloppsbanor	orbit	orbits
omnämns	is mentioned
område	area
områden	area
områdena	the areas
området	the area
områdets	the area's	of the area
omröstning	vote
omröstningen	vote	the election
omskärelse	circumcision
omslaget	cover	the cover
omstritt	controversial
omständigheter	circumstances
omtvistat	contentious	disputed	controversial
omvandlar	transmuted
omvandlas	convert
omvandling	transformation
omvända	reverse
omvänt	reversed	vice versa
omvärlden	surrounding world	outside world
omväxlande	varied
omöjligt	impossible
on	on
onani	masturbation
onda	evil
ondska	evil
ondskan	the evil	evil
ont	bad
ontario	ontario
open	open
opera	opera
operan	opera	the opera
operation	operation
operationer	operations
operativsystem	operating system	operative systems	os
opinion	opinion
opinionen	opinion
opposition	opposition
oppositionen	opposition
oralsex	oral sex
orange	orange
ord	word
ordagrant	literally	literal
ordbok	dictionary
orden	the words	words
ordentligt	proper	properly
ordet	the word	word
ordförande	chairman
ordinarie	permanent	ordinary	regular
ordna	arranging	arrange
ordnade	arranged
ordnar	fix	decorations
ordning	system
ordningen	the order	order
ordspråk	proverb	saying
organ	body	agency	organ
organisation	body	organization
organisationen	the organization
organisationens	the organizations
organisationer	organizations	organisations
organisera	organize	organizing
organiserad	organised	organized
organiserade	organized
organiseras	organizes	organized
organiserat	structured
organisk	organic
organiska	organic
organism	organism
organismen	the organism
organismer	organism	organisms
orgasm	orgasm
origin	origin
original	original	orignal
orkester	orchestra
ormar	snakes
oro	worry	concern
orolig	worried
oroligheter	unrest
orsak	reason	cause
orsaka	cause
orsakad	caused	induced
orsakade	caused
orsakar	causes
orsakas	caused	causes
orsakat	caused
orsaken	reason	cause
orsaker	causes
orsakerna	the causes
ort	neighborhood	place	location
orten	the suburb
orter	locations	varieties
ortodoxa	orthodox
os	os
oscar	oscar
oskar	oskar
oslo	oslo
osmanerna	ottoman turks
osmanska	osmanian	ottoman; osmanli
oss	center	us
ost	cheese
osv	etc.
osäker	insecure	unsure
osäkert	insecure	uncertain
osäkra	insecure
otaliga	countless; endless	countless
otto	otto
out	out
ovan	above
ovanför	over	above
ovanlig	unusual	uncommon
ovanliga	unusual	rare
ovanligt	unusual
ovanpå	on top of
ovanstående	above
oväntat	unexpectedly	unexpected
own	egen
oxenstierna	the oxenstierna
oxford	oxford
ozzy	ozzy
oändligt	infinitely
pablo	pablo
page	page
pakistan	pakistan
palats	palaces	palace
palestina	palestine
palestinier	palestinians	palestinian
palestinsk	palestinian
palestinska	palestinian
palme	palme
palmes	palme's	plame's
pamela	pamela
panthera	panthera
pappa	dad
papper	paper
par	pair
paradiset	the paradise	paradise
paraguay	paraguay
parallella	parallel
parallellt	parallel
parentes	brackets
paret	pair	the couple	parathyroid
paris	paris
park	park
parken	park	the park
parker	parker
parlament	parliament
parlamentarisk	parliamentary
parlamentariska	parliamentary	the parliamentary
parlamenten	parliaments	the parliament
parlamentet	the parlament	parliament
parlamentets	the parliament's
parlamentsvalet	parliament election	election to parliament
parten	party
parter	party
parterna	parties
parti	party
partido	partido
partier	portions	parties
partierna	portions
partiet	the party	portion
partiets	the party's	parties
partiklar	particles
partiledare	party leader
partner	partner
partnern	the partner
pass	an
passa	fit
passade	suiting	suited	fit; suited
passagerare	passenger
passagerarna	passengers	the passengers
passande	fitting	suitable	matching
passar	suits
passera	pass
passerade	passed
passerar	passes
passiv	passive
pastor	pastor
pastoral	pastoral
patent	patent
patienten	the patient
patienter	patients
patrick	patrick
patrik	patrik
patterson	patterson
paul	paul
paulo	paulo
paulus	paulus	paul
paus	pause	paus
paz	paz
pc	pc
peang	hemostat	clamp	hemostatic forceps	forceps	hemostatic clamp
pearl	pearl
peka	point (at; to; in)	point
pekar	points	pointer	pointing
pekat	pointed	identified
peking	beijing
pelle	pellet
pendeltåg	commuter train	commuter
pengar	money
pengarna	the money	money
penis	penis
pennsylvania	pennsylvania
people	people
per	per
perfekt	perfect
performance	uppträdande
period	period
perioden	period	time
perioder	periods; episodes	period
periodiska	periodic
periodvis	periodically
permanent	permanent
permanenta	permanent
pernilla	pernilla
perro	perro
perry	perry
persbrandt	persbrandt
perserna	the persians	persians
persien	persia
persiska	persian
person	person
personal	personal	employed	staff
personalen	the staff
personen	the person
personens	the persons	the person's
personer	person	people
personerna	people; persons	the persons
personlig	personal
personliga	personal
personligen	individual	personally
personlighet	character	personality
personlighetsstörning	personality disorder
personlighetsstörningar	personality disorders
personligt	personal
persons	a person's	persons	person's
perspektiv	perspective
persson	persson
peru	peru
peruanska	peruvian
pest	plague
pesten	the plague
peter	peter
peters	peters
petersburg	petersburg
petra	petra
petroleum	petroleum
petrus	petrus
petter	petter
pettersson	pettersson
pga	because of (short of "på grund av")
ph	ph
phil	phil
philadelphia	philadelphia
philip	philip
philips	philips
phoebe	phoebe
phoenix	phoenix
pi	pi
piano	piano
picasso	picasso
picchu	picchu
picture	picture
pierre	pierre
pilatus	pilatus	pilate
pink	pink
pippi	pippi
pippin	pippin
pirate	pirate
piratpartiet	pirate party
pitt	pitt
pjäs	piece
pjäsen	play
pjäser	plays
place	place
placera	position	place
placerad	placed
placerade	put	placed	placed (in)
placerades	placed
placerar	place	places
placeras	placed
placering	placement
plan	level
planen	the field	the plan	plan
planer	plans
planerad	planned
planerade	planned
planerar	is planning	plan
planeras	is planned	planned
planerat	planned
planering	planning
planerna	the plans	plans
planet	planet
planeten	the planet
planetens	planet	the planets
planeter	planets
planeterna	the planet's	the planets
planeternas	the planets'	planets	the planets
plasma	plasma
platina	platinum
platon	platon	platonic
platons	platon's	platos
plats	place	place; position
platsen	the place	place
platser	places
platt	flat	plate
platta	flat
plattan	plate	the plate
plattform	stage; platform	platform, pad, rig	platform; stand	platform, pad, stand	platform	plattform
platån	the plateau	plateau
player	player
playstation	playstation
plikt	duty
plikter	duties
plocka	pick
plural	plural
plus	plus
pluto	pluto
plötsligt	suddenly	sudden
poe	poe
poes	poe's	poes
poesi	poetry
poet	poet
poeten	poet	the poet
poeter	poets
point	point
pojkar	boys
pojkarna	boys	the boys
pojke	boy
pojkvän	boyfriend
polacker	polish	poles
polen	poland	pole
polens	polands
policy	policy
polis	police
polisen	police	the police
polisens	police	the police's
poliser	police (-men; -women)	police
politik	politics	policies
politiken	the politics
politiker	politicians	politician
politisk	political
politiska	politic
politiskt	political
polska	polish
pommern	pommern	pomerania
pompejus	pompejus
ponny	pony
pontus	pontus
pop	pop
popsångare	popsinger	pop singer
popularitet	popularity
population	population
populationen	the population	population
populationer	populations
populär	popular
populära	popular
populäraste	rated	most popular
populärkultur	popular culture	pop-culture
populärkulturen	popular culture
populärmusik	popular music	pop music
populärt	popular	popularly
port	gate
porto	postage
porträtt	portrait
portugal	portugal
portugals	portugals	portugal
portugisiska	portuguese	portugese
position	position
positionen	position	the position
positioner	positions
positiv	positive
positiva	positive
positivt	positive
post	not a swedish word
posten	the position
poster	positions	post offices
postumt	posthumously
potatis	potato
potential	potential
potentiellt	potential
potter	pots	potter
povel	povel
poäng	score	point
prag	prague
praktiken	practice	practically
praktisk	practical
praktiska	practical
praktiskt	convenient
prata	talk
pratar	talks	talking
praxis	practice
precis	precisely	exactly; precisely
premier	premiums
premiär	premiere
premiären	premiere	premier
premiärminister	prime minister
premiärministern	the prime minister	prime minister
preparat	substance	compound
presenterade	presented
presenterades	presented
presenterar	presents	present
presenteras	was presented	presented
president	president
presidenten	the president
presidentens	the president's	president	the presidents
presidenter	presidents	president
presidentvalet	presidential elections	presidential election
presley	presley
press	press
pressas	pressed
pressen	press	the pres
prestigefyllda	prestigious
preussen	prussia
preventivmedel	contraceptives
primitiva	primitive
primtal	prime number
primära	primary
prince	prince
princip	principle	principal
principen	the principal
principer	principals	principles
prins	prince
prinsen	prince	the prince
prinsessan	the princess	princess
pris	price	prize
priser	rates	prizes
priserna	prices	the prices
priset	the prize
prisma	prisma	prism
pristagare	laureate	prizewinner
privat	private
privata	private
privatliv	private
privilegier	privileges
privilegium	privilege	prerogative	privelege
problem	problem
problemen	problems	the problems
problemet	the problem
procent	percent	per
process	process
processen	process	the process
processer	processes
producent	producers	prodcuer	producent; tillverkare	producer
producenten	the producer	producer
producenter	producers
producera	produce
producerad	produced
producerade	produced
producerades	was produced
producerar	producing	produces
produceras	produced
producerat	produced
producerats	produced	produced (by)
produkt	product
produkten	product	the result
produkter	products
produktion	production
produktionen	the production
produktiv	productive
professionell	professional
professionella	professional
professor	professor
professorn	professor	the professor
profet	prophet
profeten	the prophet
profeter	prophets	profets
profil	profile
programledare	host
programmet	the application	the program
programvara	software
projekt	project
projektet	project
prokaryoter	prokaryote
promemoria	short essay	memo	memorandum	aide-memoire	pm; memorandum	promemoria
propaganda	propaganda
proportioner	proportions
prosa	prose
protein	protein
proteiner	proteins
proteinerna	the proteins	proteins
proteinet	the protein
protestanter	protestants
protestantiska	protestant	protestantic
protester	protests
protesterade	protested
protesterna	protests	the protests
protokoll	protocol
protoner	protons
prov	tests
provins	province
provinsen	the province
provinser	provinces
provinserna	the provinces
provisoriska	provisional
prägel	character	mark
präglad	characterize	characterized	marked
präglade	characterized
präglades	was marked	imprinted
präglas	characterized
präglats	marked
präster	priests
ps	ps	p.s
psykisk	psychic
psykiska	psychic	mental
psykiskt	psychic
psykologi	psychology
psykologin	the psyhology	psychology
psykologisk	psychological
psykologiska	psychological
psykos	phychosis	psychosis
psykosen	the psychosis
psykoser	psychoses
psykoterapi	psychotherapy
psykotiska	psychotic
publicera	publish
publicerad	published
publicerade	published
publicerades	published
publiceras	publishes	published
publicerat	published
publiceringen	the publication	publishing	publication
publik	audience	public
pucken	the puck
puerto	puerto	port
puls	pulse
pund	pound
punk	punk rock	punk	para
punkt	item	point
punkten	the point	point
punkter	points	seq
purple	purple
pythagoras	pythagoras
päls	fur
pär	pär
på	on	in, on, at
påbörjade	started
påbörjades	commenced; begun	initiated	was started
påbörjas	starts	start
påföljande	subsequent
pågick	lasted
pågående	current	ongoing
pågår	(in) progress
påminde	reminded
påminner	reminds	out
påsk	easter
påsken	easter
påstod	claimed
påstådda	said	alleged
påstående	assumption
påståenden	claims	assertions
påstår	claims	asserts
påstås	claimed	(been) said
påtagligt	substantially	considerably
påtryckningar	pressures	pressure
påven	the pope
påverka	influence
påverkad	influenced	affected
påverkade	influenced	affected
påverkades	was affected by	affected
påverkan	impact	influence
påverkar	affecting
påverkas	affected
påverkat	influenced
påverkats	influenced	affected
påvisa	prove	show
q	q
queen	drottning
queens	queen
rachel	rachel
rachels	rachel's
rad	range	line
radie	radius
radikala	radical
radikalt	radical	radically
radio	radio
radioaktiva	radioactive
radioaktivt	radioactive
radion	the radio	radio
rafael	rafel
ragnar	ragnar
raid	raid
rainbow	rainbow
rak	straight	linear
raka	straight
rakt	straight
ramadan	ramadan
ramel	ramel
ramels	ramel's
ramen	frame
rammstein	rammstein
rankas	ranks
rankning	ranking	rating
rankningar	rankings	ranking
rapport	report
rapporten	report	the report
rapporter	reports
rapporterade	reported
rapporterar	reports
ras	race
rasade	collapsed
rasen	breed	the race
raser	species
rasism	racism
rastafari	rastafarian
rastafarianer	the rastafarian	rastafarian	rastafarians
rastafarianerna	the rastafarian	rest are faria
reagan	reagan
reagans	reagan's
reagera	reacting
reagerar	reacts
reaktion	reaction
reaktionen	reaction	the reaction
reaktioner	reactions
reaktionerna	the reactions	reactions
reaktorer	reactors
reaktorn	the reactor	reactor
realiteten	de facto	reality
rebecca	rebecca
recensioner	reviews
receptorer	receptors
red	eds
reda	find out	out	find our
redaktör	editor
redan	already	has already
rede	clutch	nest	coated
rederiet	the shipping company	the company	shipping company
redo	ready
redovisas	shown	accounted for
redskap	device
reducera	reduce
reduktion	reduction
referens	reference
referenser	references
refererar	refer (to)
reform	reform
reformationen	the reformation
reformer	reformers	reforms
regel	rule
regelbunden	regular
regelbundet	regularly	regularily
regelbundna	regular
regeln	the rule	rule
regent	ruler	regent
regenter	monarchs
regerade	reigned
regerande	ruling
regering	the government	government
regeringar	governments
regeringen	the government	government
regeringens	government
regeringschef	head of government	government
regeringsmakten	govermental power	government power
regeringstid	term of government	term of government; term of office
reggae	reggae
reggaen	reggae	the reggae
regi	direction
regim	regime
regimen	regime
regimer	regimes
region	region
regional	regional
regionala	regional
regionalt	regional	regionally
regionen	the region
regioner	regions
regionerna	regions
regisserad	produced	directed
regissör	director
regissören	director
registrerade	data	noted
regler	rules
reglera	controlling	expell
reglerar	regulates
regleras	is regulated	regulated
reglerna	rules	rules; regulations
regn	rain
regnar	rains	raining
regnskog	rain forest	rainforest
reguljära	regular
reidar	reidar
reidars	reidar's	reidars
reinfeldt	reinfeld	reinfeldt
reklam	advertising	advertisement
reklamen	the commercial	commercial; ad; advertisment
rekord	record
rekordet	the record
relaterade	related
relation	relation
relationen	the relation	ratio
relationer	relations
relationerna	the relationships	relations
relativa	relative
relativt	relatively
releasedatum	release date
religion	religion
religionen	the religion
religionens	religion's
religioner	religions
religionerna	religions	the religions
religionsfrihet	freedom of religion	religious freedom
religiös	religious
religiösa	religious
religiöst	religious
remmer	remmer
ren	deer	clean
rena	pure
rent	true	clean
renässans	renaissance
renässansen	the renaissance	renaissance
rené	rene	rené
reologi	rheology	reology
reportrar	reporters
representant	representative
representanter	representatives
representanthuset	house of representatives
representation	representation
representativ	representative
representera	represents	represent
representerade	represented
representerar	represents
representeras	represented
reptiler	reptiles
republik	republic
republika	republic
republikanska	republican
republiken	the republic of	the republic
republikens	republic's
republiker	republics
resa	travel
resan	the trip
resande	travelling
research	research
reser	travels	rise	rises
residensstad	city of residence	county seat
resolution	resolution
resor	travels	travel
respekt	respected	respect
respektive	respective
rest	remain	rest
restaurang	restaurang	restaurant
restauranger	restaurant	restaurants
reste	moved	travelled	stood
resten	the rest
rester	remains
resterande	remaining
resultat	result	results
resultaten	the results	results
resultatet	the result	result
resultera	result
resulterade	resulted
resulterar	result	results
resulterat	resulted	resulted in
resurs	resource	resources
resurser	resources
retorik	rhetoric
retoriken	rhetoric
retoriska	rhetorical
revir	territory
revolution	revolution
revolutionen	the revolution	revolution
revolutionens	revolution	the revolutions
revolutionär	revolutionary	revolutions
revolutionära	revolutionary
revs	was demolished
reza	reza
rhen	the rhine
rice	rice
richard	richard
richards	richards
richmond	richmond
rico	rico
riddare	knight
rik	rich	rish
rika	rich
rikare	richer
rikaste	the richest	richest
rike	kingdom
rikedom	riches	wealth
riken	the kingdoms	kingdoms
riket	kingdom	the land
rikets	its	the realms
riksdag	parliament; diet	the parliament
riksdagen	the parliament
riksdagens	the parliament's	the parliaments
riksdagsvalet	parliamentary election	election to parliament	parliamentary elections
riksförbundet	national association
rikskansler	chancellor
riksrådet	privy council; council of state; crown council; senate	privy council
riksväg	national highway	highway
rikt	target	rich
riktad	directed
riktade	targeted
riktar	target	targets
riktas	directed (at)	direct
riktat	pointed
riktig	real
riktiga	real
riktigt	real
riktlinjer	guidelines
riktning	direction
riktningar	directions	direction (-s)
riktningen	direction	denomination
ring	ring
ringa	call
ringar	rings
ringde	called
ringen	ring
rinner	running	flow
ris	rice
risk	risk
risken	the risk	risk
risker	risks
riskerar	risks
rita	paint	draw
ritualer	rituals
rivalitet	rivality	rivalry
river	river
rna	rna
rob	rob
robbie	bobbie	robbie
robert	robert
roberto	roberto
roberts	roberts
robin	robin
robinson	robinson
rockband	rock band
rocken	the rock	rock
rockgrupper	rock groups	rock bands
rocksångare	rock singers	rock singer
rod	rod
roger	roger
roland	roland
roll	role
rollen	role	the role
roller	roles
rollfigur	character
rollfigurer	roll model	role figure
rolling	rolling
rom	rome	rom
roma	roma
roman	novel
romance	romance
romanen	novel
romaner	novels
romani	romany	roma
romantiken	romance	romanticism
romantikens	the romanticism	romantick
romantiska	romantic
romarna	the roman	the romans
romarriket	the roman empire
romeo	romeo
romer	romani people	roma
romerna	roma	the romani	the romani people
romersk	roman
romerska	roman
romerske	roman
romerskkatolska	roman catholic
roms	rome's	romes
romska	romani
romulus	romulus
ron	ron
ronaldinho	ronaldinho
ronaldo	ronaldo
ronden	round
ronja	ronja
roosevelt	roosevelt
rorsman	helms man	helmsman	steersman
rosa	pink	rosa
rose	rose
rosenberg	rosenberg
rotation	rotation
roterande	rotating
roterar	rotates
rousseau	rousseau
rovdjur	predator	predators
rowling	rowling
roy	roy
rubiks	rubik's
rubrik	headline	header	head line; rubric	heading	title
rudolf	rudolf
rugby	american fotboll	rugby
ruiner	ruins
rum	(took) place
rummet	room
rumänien	romania
rumänska	romanian
run	run
runda	round
running	running
runor	runes
runorna	the runes
runstenar	runestones	rune stones
runt	around	between
runtom	throughout	around
ruset	the fuddle
rush	rush
russell	russell	rusell
rwanda	rwanda
ryan	ryan
rybak	rybak
rygg	back	dorsal
ryggen	the back
rykte	reputation
rykten	rumors
rymden	space
rymmer	has	holds
rysk	russian
ryska	russian
ryssland	russia
rysslands	russia's
rytmiska	rhythmic
räcker	enough
räckte	enough	handed
rädd	scared	afraid
rädda	save	lot of
räddade	saved
räddar	saves	saved
rädsla	fear
räkna	count
räknade	calculated	counted
räknar	counts
räknas	calculated	counted	are counted
räknat	calculated	counted
rätt	right
rätta	correct	come to grips; court; correct
rättegång	trial	steering wheel gang
rättegången	trial	the trial
rätten	the court
rätter	dishes
rättigheter	rights
rättigheterna	the rights	rights
rättsliga	justice	legal
rättvisa	justice
råd	advice	council
rådande	current	prevalent
rådde	prevailed	was
råder	advises	(that) prevails
rådet	the council	council
rådets	council
rådgivare	counsellor	advisor
rådhus	courthouse
råkar	happens	happens to
råolja	crude oil
råvaror	raw	wood	raw materials
röd	red
röda	red
röka	smoke
rökning	smoking
rör	touch, move(-s)	touches	row
röra	move
rörande	concerning
rörde	had something to do with	touched	was about
rörelse	movement
rörelsen	movement
rörelsens	movement	movements
rörelser	movements
rörelserna	the movements
rörlighet	movement
röst	voice
rösta	vote
röstade	voted
rösten	the voice	rust
röster	votes
rösterna	votes	the votes
rösträtt	right to vote
rött	red
rötter	roots
sa	said
saab	saab
sabbath	sabbath
sachsen	sachsen	saxony
saddam	saddam
sade	said
sades	said	was said
saga	saga	story
sagan	story
sagor	fairytales	tales	fairy tales
sagt	said
sahara	sahara
sahlin	sahlin
saint	saint
sak	thing	matter; case
saken	the thing	the matter
saker	things
saknade	lacked	missed
saknades	lacked	missing
saknar	lacks	lack(-s)	missing
saknas	missing
sakrament	sacrament
sakta	slowly
salt	salt
salvador	salvador
sam	co
samarbeta	collaborate	cooperate
samarbetade	collaborated	collaboration
samarbetar	cooperates	collaborates
samarbetat	collaborated	collobrated
samarbete	collaboration
samarbeten	collaborations	cooperations
samarbetet	co	the collaboration
samband	connection
sambandet	the connection	connection	relation
same	lapp	sami
samerna	the lapp
samfund	communities	order
samfundet	the communion	association
samhälle	society
samhällen	communities	societies
samhället	the society	society
samhällets	society	of society
samisk	samian	lapp
samiska	sami
samla	collect	gather
samlade	collected
samlades	collected	gathered	were united
samlag	intercourse
samlar	collect	collectors
samlat	gathered
samlats	gathered; collected
samling	concentration	collection
samlingar	collections	collection
samlingsalbum	compilations
samma	the same	same
samman	together
sammanfaller	coincides
sammanfattning	summary
sammanhang	context
sammanhanget	connection	context
sammanhängande	continous	connective
sammanlagt	a total of
sammansatt	composed
sammansatta	composed	joined
sammansättning	composition
samoa	samoa
samspel	interaction	teamwork
samt	also	as well as
samtal	call	conersation
samtida	contemporary
samtidigt	while	simultaneous
samtliga	all
samtycke	approval
samuel	samuel
samverkan	co	cooperation
samverkar	co-operating	co-operates
samväldet	commonwealth	the commonwealth
san	san
sand	sand	sandy
sandy	sandy
sankt	sankt	st.
sankta	sankta	saint
sann	true
sanna	true
sanning	truth
sanningen	the truth
sannolikhet	probability
sannolikt	probable
sanskrit	sanskrit
sant	true
santa	santa
santiago	santiago
sapiens	sapiens
sara	sara
sarah	sarah
sarajevo	sarajevo
satan	satan
satanism	satanism	satanic
sats	statements	clause	sets	kit	proposition	statement	theorem	theorems; sets	proof	theorem; sets
satsa	bet
satsade	bet
satsningar	investments	resources
satt	saat	sat
satte	put	put together	sat
sattes	was added
saturnus	saturnus
saudiarabien	saudi arabia
sauron	sauron
sawyer	sawyer
scen	scene
scenen	the stage
scener	scenes
schack	shack	schack	chess
schizofreni	schizophrenia
schwarzenegger	schwarzenegger
schweiz	switzerland
schweiziska	swiss
science	science
scientologikyrkan	the church of scientology	church of scientology
scott	scott
screen	screen
se	see
sean	seab	sean
sebastian	sebastian
sed	thirst
sedan	then	since
sedd	seen
seden	the seed	custom
seder	custom
sedermera	subsequently	since
sedlar	bills
seger	victory
segern	the victory	victory
seglade	sailed
segrar	wins	victories
sekel	century
sekelskiftet	turn	the turn of the century
sekreterare	secretary
sekt	sect
sekter	sects
sektion	section
sektorn	sector	the sector
sekulär	secular
sekulära	secular
sekunder	seconds	second
sekvens	sequence
selassie	selassie
selma	selma
semifinal	semi finals
semifinalen	semi finals
sen	then	since
sena	late
senare	latterly; later	later
senast	last (time)	last
senaste	last
senaten	senate	the senate
senator	senator
sent	late
sentida	recent
separat	seperate	separate
separata	separate
separerade	separated
september	september
ser	see	sees
serber	serbs
serbien	serbia
serbiens	serbias
serbisk	serbian
serbiska	serbian
serie	comic; row; succession; serial	cartoon	series
serien	the series
seriens	series
serier	comics
serotonin	serotonin
serveras	is served
service	service
servrar	servers
ses	are seen
seth	seth
sett	seen
setts	seen
sevärdheter	attractions
sex	six
sexton	sixteen
sexualitet	sexuality
sexuell	sexual
sexuella	sexual
sexuellt	sexual
sfären	sphere
shahen	the shah	shah
shakespeare	shakespeare
shakespeares	shakespeare's
sharia	sharia
sheen	sheen
sibirien	siberia
sicilien	sicily
sida	website	side
sidan	page	the side	side
side	side
sidor	pages
sidorna	the pages	pages
sierra	sierra
siffra	number
siffran	number	the number
siffror	numbers
siffrorna	the numbers	numbers
sig	to	itself
sigmund	sigmund
signaler	signals
signifikant	significant
sikt	run
silver	silver
simmons	simmons
simning	swimming
simon	simon
simpson	simpson
simpsons	simpsons
sin	its
sina	their
sinatra	sinatra
singapore	singapore
singapores	singapores	singapore's
singel	single
singeln	single
singer	singer
singlar	singles
singlarna	the singles
sinne	mind
sir	sir
sist	last
sista	last
siste	lattermost	last
sistnämnda	later
site	site
sitt	his	its
sitta	sit
sittande	fitting	sitting
sitter	serve	sit
situation	situation
situationen	situation	the situation
situationer	situations
siv	siv
sixx	sixx
sju	seven
sjuk	ill	disease
sjuka	disease	sick
sjukdom	illness	disease
sjukdomar	diseases	disease
sjukhus	hospital
sjukhuset	the hospital	hospital
sjukvård	health care	care	healthcare
sjunde	seventh
sjunga	access	sing
sjunger	sings	singing
sjunka	decrease	descend
sjunkande	sinking; decreasing	decreasing
sjunker	sinks
sjunkit	decreased
själ	soul
själen	the soul
själv	own	alone	himself
själva	self	actual
självbiografi	autobiography	selfbiografi
självklart	course
självmord	self-killing	suicide
självstyrande	independent	self-governance
självstyre	autonomy	self-governance
självständig	independent	independant
självständiga	independent	sjalvstandiga
självständighet	independance	independence
självständigheten	independance	independence
självständigt	independent	independant
självt	itself
sjätte	sixth
sjö	lake	naval
sjöar	lakes	parks
sjöarna	the lakes	lakes
sjöfart	sea voyage	navigation
sjöfarten	shipping
sjögren	sjögren
sjön	lake
sjöng	sang
sjönk	decreased	sank	sunk
sjöss	sea
sk	so called	known
ska	will
skabb	scab	scabies
skada	damage
skadad	damaged
skadade	wounded	damaged
skadades	was wounded
skadan	damage	the damage	the hit
skadas	damaged
skadliga	harmful	deleterious
skador	damage
skadorna	damages	injuries	damage
skaffa	obtain	gain
skaffade	aquired
skal	shell
skala	scale	scale; size
skalan	scale
skalet	shell	the shell
skall	is	shall
skalv	quake
skalvet	quake
skandinavien	scandinavia
skandinaviska	scandinavic	scandinavian
skapa	create
skapad	created
skapade	made	created
skapades	created
skapande	building	creating	creative
skapandet	creation	the making
skapar	creates
skapare	creator
skapas	creates
skapat	created
skapats	was created	generated
skapelse	creation
skara	city in south-central sweden (uppland)
skarp	sharp	crisp
skarsgård	skarsgård
skatt	tax
skatter	taxes
ske	be	happen
skedde	was
skede	period
skelett	skeleton
skepp	ship
skeppen	the ships
skeppet	the ship
sker	happens	is
skett	happened
skick	state
skicka	send
skickade	sent
skickades	was sent	sent
skickar	sends	send
skickas	is sent
skicklig	skillful	proficient	skilled; skillful
skiftande	shifting
skikt	layers
skilda	seperated	separate
skilde	divided
skildes	separated	was seperated
skildrar	describes	portrays
skildras	is depicted
skildringar	description	descriptions
skilja	seperate	differ; differentiate	separate
skiljas	separate
skiljer	differs	is different; differ
skiljs	separated	separate
skillnad	difference
skillnaden	the difference
skillnader	differences
skillnaderna	the differences
skilsmässa	divorce
skiva	record	disc
skivan	record	the record	disc
skivbolag	record label	record company
skivbolaget	record label	the record company
skivkontrakt	record deal	record contract
skivor	plates	records
skivorna	the records	records	plates
skjuta	delay	postpone; shoot
skjuten	shot
skjuter	shoots
skog	wood	forest
skogar	forests
skogarna	the forests	forests
skogen	woods	forest
skola	school
skolan	school
skolgång	school attendance	schooling
skolor	schools
skolorna	the schools
skor	shoes
skorpan	crust
skotsk	scottish
skotska	scotland	scottish
skott	round	shots
skottland	scotland
skov	episode	relapse
skrev	said
skrevs	written	was
skrift	book	writing
skriften	no.	writings
skrifter	writings
skrifterna	scriptures
skriftliga	written
skriva	write
skrivas	written
skriven	written
skriver	write	type
skrivet	written
skrivit	written	wrote
skrivits	been written
skrivna	written
skrivs	written	printed
skräck	horror	fear
skuggan	the shadow
skuld	debt	guilt
skulden	the debt	the guilt
skulder	liabilities	debts	debt
skull	sake
skulle	could	would
skulptur	sculpture
sky	sky
skydd	protection
skydda	protect
skyddade	protected
skyddar	protection	protects
skyddas	(is/are) protected
skyldig	responsible	guilty
skyskrapor	high rise buildings; sky scrapers
skäl	reasons	reason
skär	will	skerry
skära	carve	cut
skärgård	archipelago	archipelagos
skådespelare	actor
skådespelaren	actor
skådespelarna	actors
skådespelerska	actress
skåne	skåne
skånes	scania's
skånska	scanian dialect	scanian	skånska
skönhet	beauty
skönlitteratur	fiction
sköt	shot
sköta	operate	handle
sköter	handles	handle
sköts	postponed; run	shot	handled
sköttes	operated	handled
slag	type	kinds
slaget	the strike
slagit	held	beaten
slags	kind	type
slavar	slaves
slaveriet	slavery
slaviska	slav	slavic
slidan	the vagina	vagina
slipknot	slipknot
slippa	avoid
slog	hit
slogs	fought	was
slott	castle
slottet	the castle
slovakien	slovakia
slovenien	slovenia	slovenian
slovenska	slovenian
slut	end
sluta	end
slutade	quit
slutar	ends	end
slutat	ended
slutet	end
slutgiltiga	final
slutliga	evenutal	ultimate
slutligen	at last
slutsats	conclusion
slutsatsen	the conclusion
slutsatser	conclusions
släkt	family
släkten	the family
släktet	the genus
släkting	relative
släktingar	relatives
släktskap	relationship	kinship
släppa	release
släppas	released	be released
släpper	release	releases
släpps	released	(is) released
släppt	self-indulgent	released	relinquished
släppte	released
släpptes	was released
släppts	released
slå	hit
slår	states	beats
slås	beat	is hit	slas
slåss	fight
slöt	joined (in peace)	closed
slöts	concluded	signed
sm	s-m	swedish championship
smak	taste
smaken	the flavour	flavor
smala	narrow
smallwood	small wood	smallwood
smeknamn	nickname
smeknamnet	nickname
smguld	swedish championship gold	gold medal in the swedish championships
smith	smith
smitta	infection
smycken	jewlery
smält	melted
smärta	pain
små	little, small	small
småland	smaland
smålands	smaland's
småningom	eventually
snabb	instant
snabba	rapid	fast
snabbare	rapid	faster
snabbast	fastest
snabbaste	rapid	fastest
snabbt	quickly
snarare	rather
snarast	rather	as soon as possible
snart	soon
snitt	on average	average
snittet	average
snus	snuff
snuset	snuff	the snuff
snö	snow
social	social
sociala	social
socialdemokrater	social democrats
socialdemokraterna	members of the social democracy
socialdemokratiska	socialists	social democratic
socialism	socialism
socialismen	the socialism	socialism
socialister	socialists
socialistisk	socialistic	socialist
socialistiska	socialistic
socialistiskt	socialistic	socialist
socialt	social
socken	parish
socker	sugar
sofia	sofia
sofie	sofie
sokrates	socrates	sokrates
sol	sun
soldat	soldier
soldater	soldiers
soldaterna	soldiers	the soldiers
solen	the sun	sol
solens	the sun
solljus	sun light	sunlight
soloalbum	solo album
solsystem	solar system
solsystemet	the solar system	solar system`
solsystemets	solar system
solvinden	the solar wind
som	as	which
somalia	somalia
somliga	some
sommar	summer
sommaren	the summer
sommarspelen	summer games
sommartid	summer-time	during summer
somrar	summers
somrarna	the summers	summers
son	son
sonen	the son
sony	sony
sorg	grief
sorter	kinds	types
sorters	kinds	kinds of
sorts	variety
soul	soul
sound	sound
soundtrack	soundtrack
south	south
sover	sleep
sovjet	soviet
sovjetisk	soviet	sovietic
sovjetiska	soviet	sovjet
sovjetunionen	the soviet union
sovjetunionens	soviet union's; soviet's	soviet union
spaniel	spaniel
spanien	spain
spaniens	spain's
spanjorerna	the spaniards	spanish
spannmål	cereals	grain
spansk	spanish
spanska	spanish
sparken	park	fired	gets fired
sparta	sparta
spears	spears
special	special
specialiserade	specialized
speciell	special
speciella	special
specifik	specific
specifika	specific
specifikt	specifically
speglar	mirror	mirrors
spektrum	spectra	spectrum
spektrumet	spectrum
spekulationer	speculations
spel	game
spela	play
spelad	played
spelade	played
spelades	filmed
spelar	gaming
spelare	player
spelaren	the player
spelarna	players
spelas	played
spelat	played
spelats	been played	played
spelen	the games
spelet	the game
spelfilmer	motion pictures	feature film	feature films
spelning	gig	playing
spelningar	tour	gigs
spelningen	the gig
spets	edge; top	point
spetsen	edge; top
spetshundar	tip of dogs
spindlar	spiders
spindlingar	slindlingar	cortinariuses	webcap	spindlingar	fungus	cortinarus	spiders	cortinarius	cortinariaceae	this is not a swedish word.
splittrades	shattered	split
spontant	spontaneous	spontaneously
sport	athletics	sport
sporten	the sport
sporter	sports
spotify	spotify
spred	spread
spreds	spread	disseminated
sprida	spread
spridas	spread
spridd	spread
spridda	spread	scattered
sprider	spreads out	spread	spreads
spridit	spread
spridning	diffusion	distribution
spridningen	spread	the spread
sprids	spreading	spreads
springer	running
springsteen	springsteen
springsteens	springsteen's	springsteens
sprit	liqeur	alcohol
spritt	spread
språk	language
språkbruk	parlance	language (use); parlance; phraseology
språken	languages	park
språket	language
språkets	the language's	language
språkliga	linguistic
spänner	span
spänning	voltage
spänningar	tensions
spänningen	exitement	voltage
spår	track	pairs
spåra	track	trace
spåras	trace
spåren	the tracks	tracks	wake
spårvagnar	trams
sr	sr
sri	sri
ss	ss
st	saint
stabil	stable
stabila	stable
stabilitet	stability
stad	city
staden	the city
stadens	the town's	the citys	city's
stadigt	stable	steadily
stadion	stadium	the stadium
stadium	stage
stadsbild	cityscape
stadsdel	city district	district
stadsdelar	districts	city districts
stadsdelarna	districts	neighborhood (-s)
stadsdelen	the district
stadshus	city hall; town hall	town hall
stadskärna	city core, city center	town centre
stadskärnan	town/city	center
stadsparken	city park	city ​​park
staffan	staffan
stalin	stalin
stalins	stalins	stalin
stallone	stallone
stam	tribe
stammar	tribes	stutters
stammarna	tribes
stan	town
stand	stand
standard	standard
stanley	stanley
stanna	stay
stannade	stayed
stannar	stays	stop	stay
stark	strong
starka	strong
starkare	strong	stronger
starkast	strongest
starkaste	strongest	the strongest
starkt	strongly
start	start
starta	launch
startade	started
startades	started
startar	begins	starts
startat	started
starten	the start	start
stat	state
state	state
statens	state	the government's
stater	states
staterna	usa
staternas	states	the state's
states	states
station	station
stationen	station
stationer	stations
statistik	statistics
statistiska	statistical
statlig	state	government
statliga	state
statligt	governmental
stats	state's
statschef	head of state
statschefen	the head of state	head of state
statskupp	coup
statsmakten	the government	power	government
statsminister	prime minister
statsministern	prime minister	head of state
statsreligion	state religion
statsskick	polity	form of government
statsöverhuvud	head of state
status	status
staty	statue
statyn	the statue
stavning	spelling
stavningen	spelling	the spelling
stefan	stefan
steg	rose	step
steget	step
sten	stone
stenar	stones	blocks
stephen	stephen
steve	steve
steven	steven
stewart	stewart
stieg	stieg
stift	pin	diocese
stiftelsen	foundation
stig	stig
stiga	rise
stigande	rising
stiger	rises
stilar	styles
stilen	style
stilla	still
stimulans	stimulation	stimulating
stimulera	stimulate	stimulating
stimulerar	stimulates
stjäla	steal
stjärna	star
stjärnan	star	the star
stjärnans	star's	the star's	the stars
stjärnor	stars
stjärnornas	the star's
stockholm	stocholm	stockholm
stockholms	stockholm's	stockholm
stod	stood
stoft	dust
stol	chair
stolpiller	suppository	pauropoda	stolpills	suppositary
stommen	frame	the foundation
stop	stop
stopp	stop
stoppa	stop
stoppade	stop	stopped
stor	big; great
stora	large	big
storbritannien	great britain	uk
storbritanniens	uk
store	great
stores	the great	the great's
storhetstid	heyday
storkors	the grand cross
storlek	size
storleken	size
storm	storm
stormakt	great power
stormakter	world powers	great power	superpowers
stormakterna	great powers
stormaktstiden	great power period	greatness
storstäder	metropolises	cities
stort	large	big
stortorget	stortorget	the main square
story	story
straff	punishment	punishments
straffet	penalty	the punishment
strand	beach
stranden	shore	the beach
strategiska	strategical	strategic
stratton	stratton
strax	soon	just
streck	bar
stred	fought
street	street
stress	stress
stressorer	stressors
strid	fight
strida	fight
stridande	fighting
striden	fight
strider	conflict	battles
striderna	the battles	fighting
stridigheter	oppositions
strikt	strict
strikta	strict
strindberg	strindberg
strindbergs	strindberg's
struktur	structure
strukturen	the structure
strukturer	structures
sträckan	the distance
sträcker	stretches	extend
sträckor	distances
sträckte	extended
stränder	beaches
sträng	string	strang
stränga	severe
strävan	endeavor	the quest
strävar	striving; aiming (to; for)	strives
strävhårig	hispid	wirehaired
strålning	radiation
strålningen	the radiation	radiation
ström	stream	icon
strömmar	flow	streams
strömmen	the stream
strömning	flow
strömningar	sentiments	tendencies
stuart	stuart
student	student
studenter	students
studenterna	students	the students
studera	study
studerade	studied
studerar	study	studies
studeras	(is) studied	is studied
studerat	studied
studie	study
studien	study	the study
studier	studies
studierna	studies	the studies
studiet	the study
studio	studio
studioalbum	studio album
studioalbumet	studio album
studion	studio	the studio
studios	the studio's
stulna	stolen
stund	while	momentum
stundom	sometimes	somtimes
stupade	fallen	killed
sture	sture
stycke	piece	piece; part; section
stycken	pieces; parts
styr	controls
styra	controlling	steer
styrande	rulers
styras	steered
styrde	steered
styrdes	governed	ruled
styre	rule
styrelse	government; direction	board of directors
styrelsen	the board	board
styrelseskick	form of government	government
styret	gate
styrka	strength	power
styrkan	strength; unit; force	strength
styrkor	strenghts
styrkorna	forces
styrs	is controlled	ruled
städer	urban	cities
städerna	the towns
ställa	make	set	installation
ställas	set	be set
ställde	stood up	asked
ställdes	prepared
ställe	stalle	place
ställen	spots; places	places
ställer	running; causing	run (in election)
stället	the place	instead
ställning	position
ställningar	positions	standings	notions
ställningen	position
ställs	is
ställt	put	taken	set
stämma	sue
stämmer	(if it's) true	correct
ständerna	the cities
ständig	constant
ständiga	permanent
ständigt	always	constant
stänga	close
stängdes	closed
stängt	closed
stärka	strengthen; bolster
stärkelse	starch
stärkte	strengthened	increased
stärktes	was strengthened	was strenghten
stätta	tile	start	stile	stiles
stå	stand
stående	standing
stål	steel
stålgemenskapen	steel community
stånd	in the context: (make) the war happen
ståndpunkt	standpoint
står	standing	star	stand
stått	stood
stöd	support
stödde	supported
stöder	supporting	supports
stödet	support	the support
stödja	support
stödjer	support	supports
stöds	supported	stood	is supported
störningar	interruptions	disorder	disorders
större	bigger
störst	most
största	biggest	largest
störta	rush	crash
störtades	overthrew	overthrown	was overthrown
stöter	thrust	run
stött	met
stövare	beagle	hound
substantiv	noun
successivt	successively	progressively
succé	succes	success
sudan	sudan
sugga	soe	barrier	sow
sultanen	sultan
summa	sum	total
summan	sum	the sum
summer	sommar
sun	sun
sund	sane	narrow
sundsvall	sundsvall
sundsvalls	(city of) sundsvall's
super	super
supportrar	supporters
sur	acidic	sour
susan	susan
sushi	sushi
sutra	sutra
suttit	sat
suverän	terrific	supreme	sovereign
suveräna	terrific	supreme	sovereign
suveränitet	sovereignty
sv	south west
svag	weak
svaga	faint	weak
svagare	weaker	weak
svagt	weak
svar	answer	response
svarade	accounted (for); answered	answered
svarar	responds
svart	black
svarta	black
svartån	svartån
svavel	sulphur
svealand	svealand
sven	sven
svensk	swedish
svenska	swedish
svenskan	swedish	the swede
svenskans	the swedish language	swedish language
svenskar	swedish
svenskarna	the swedes
svenske	swedish
svenskspråkiga	swedish speaking	swedish-speaking
svenskt	swedish
svensson	svensson
sverige	sweden
sverigedemokraterna	sweden democrats
sveriges	swedens	sweden
svt	svt
svält	starvation	starvations
svärd	sword
svår	severe	difficult
svåra	answering	difficult
svårare	harder
svårigheter	difficulties	hardships
svårt	difficult
swahili	swahili	swahilli
swan	swan
sweden	sweden
swedish	swedish
sweet	söt
swift	swift
syd	south
sydafrika	south africa
sydafrikanska	south african	african
sydafrikas	of south africa	south africa's
sydamerika	south america
sydeuropa	south europe	southern europe
sydkorea	south korea
sydliga	southern
sydligaste	southernmost	most southern
sydost	south east
sydostasien	south east asia
sydstaterna	the southern states	southern united states
sydväst	southwest
sydvästra	southwest
sydöst	south east
sydöstra	south east	the southeast	south eastern
syfta	aim	refer
syftade	alluded to
syftar	refers	seek to	refer
syfte	purpose
syften	purpose
syftet	purpose
symbol	symbol
symbolen	the symbol
symboler	symbols
symboliserar	symbolized	symbolizes
symbolisk	symbolic
symptom	symptoms
symptomen	symptoms	the symptoms
symtom	symptoms	symptom
symtomen	symptoms	the symptoms
syn	sight	view
synd	sin
synder	sins
syndrom	syndrom
synen	the view	sight
synes	seems to	apparently	appears
synliga	visible
synligt	visible	seen
synnerhet	specially	particular
synnerligen	remarkably; particularly	quite
synonymt	synonymous	synonymously
syns	seen
synsätt	viewpoint
synsättet	approach	view
syntes	synthesis
synvinkel	perspective
syre	oxygen
syret	the oxygen	oxygen
syrgas	oxygen
syrien	syria
syskon	sibling	siblings
sysselsätter	employs
system	system
systematik	systematic
systematiska	systematic	systematical
systematiskt	systematic
systemet	the system
systems	system	systems
syster	sister
systrar	sisters
säga	say
sägas	is said	is said (to be)
säger	says	claims; says
sägs	said (to be)	said
säker	items
säkerhet	safety; security	security
säkerheten	the security	safety
säkerhetspolitik	safety policy	security policy
säkerhetsråd	security council
säkerhetsrådet	security
säkert	securely
säkra	reliable	safe	secure
sälja	sell
säljande	selling
säljas	is sold	sold
säljer	sells
säljs	sold
sällan	seldom	rare
sällskap	company
sällskapet	the company
sällskapshundar	pet dogs	companion dog
sällsynt	rare
sällsynta	rare
sämre	poor
sämsta	worst
sända	broadcast	transmitting
sändas	broadcast	be transmitted
sände	sent
sändebud	messenger
sänder	broadcast	transmits
sändes	was sent	sent
sänds	sends	sands
sänka	lower
sänker	lowers	sinks
sänktes	sunk	reduced
särdrag	feature	features
särskild	specific	particular
särskilda	specific	special
särskilt	particulary	especially
säsong	season
säsongen	season
säsongens	season	the seasons
säsonger	seasons
säsongerna	seasons
säte	sate	seat
sätt	manner	way
sätta	insert
sättas	turn
sätter	place	puts	sets
sättet	manner	way	the way
sätts	turned (on)	is placed
så	so
sådan	such	kind of
sådana	such
sådant	such
såg	saw
sågs	seen	was observed
sålda	sold	salda
sålde	sold
såldes	sold
således	hence	thus
sålt	sold
sålts	sold
sålunda	thus
sång	song
sångare	singer
sångaren	the singer
sången	the song	song
sånger	songs
sångerna	song are	the songs
sångerska	songstress	singer
sår	sir	wound
såsom	like
såväl	both	as well as
söder	south
söderut	south
södra	southern	south
söka	search	searching
söker	searches	seeks out
sökt	searched
sökte	searched
sömn	sleep
söndagen	sunday
sönder	broken
söner	sons
t	t	e.g.
ta	to	take
tabell	table	chart	tabel
tabellen	the chart	table; list
tacitus	tacitus
tack	thanks
tackade	thanked	said/thanked
tag	while
tagen	taken
taget	a time (practically; virtually; any; at all)
taggar	spikes	thorn, twig
tagit	taken	received
tagits	taken
taiwan	taiwan
taket	the roof
takt	rate
taktik	tactics	tactic	strategy
tala	speak
talade	spoken
talades	spoken	spoken (of)	spoke
talang	talent
talanger	talents
talar	speaks	speak
talare	speaker	spoke
talas	spoken	is spoken
talat	spoken	spoke
talen	years
talet	rate	century
talets	the speechs
talman	spokesperson	speaker
talmannen	speaker of the riksdag
talrika	numerous
tankar	thoughts
tanke	light	in light of
tanken	the thought	idea
tanzania	tanzania
tappade	lost
tappar	drop	lose
tar	takes
tas	is taken
taube	taube
taubes	taubes
taylor	taylor
te	tea
team	team
teater	theatre; theater	theater
teatern	the theater	theater
teatrar	theaters
tecken	signs	sign
tecknade	cartoon (-s)	drew
tecknet	the sign	sign
ted	ted
teddy	teddy
tegel	brick
teknik	technique	technic
tekniken	techinque	the technology
tekniker	technician
teknisk	technical
tekniska	technical
tekniskt	technical
teknologi	technology
telefon	telephone
telefonen	phone	the telephone
telegram	telegram
television	television
tema	theme
teman	themes
tempel	temple
temperatur	temperature
temperaturen	temperature
temperaturer	temperature
tempererat	temperate	tempered
templet	the temple	temple
tendens	tendency
tendenser	tendencies
tenderar	tend
tenn	tin
tennessee	tennessee
tennis	tennis
tennisspelare	tennis player
teologi	teology	theology
teologiska	theological
teoretiker	theorists
teoretisk	theoretical
teoretiska	theoretical
teoretiskt	theoretic	theoretical
teori	theory
teorier	theories
teorin	the theory
termen	the term	term
termer	term
terminologi	terminology
terrier	terriers	terrier
territoriella	territorial
territorier	territories
territorierna	territories
territoriet	territory
territorium	territory
terror	terror
terrorism	terrorism
terrorismen	terrorism	the terrorism
terrorister	terrorists
terry	terry
terräng	off	terrain
tesla	tesla
teslas	tesla's
test	test
testamente	will
testamentet	testament
tex	for example
texas	texas
text	text
texten	the text
texter	texts
texterna	text
th	th
thailand	thailand
than	than
that	that
thc	thc
the	the
theodor	theodor
theta	theta
they	they
thierry	thierry
thomas	thomas
thriller	thriller
thåström	thåström	thastrom
tibet	tibet
tid	time
tiden	the time	time
tidens	time's	time
tider	times; ages	times
tiderna	the times	times, ages	time
tiders	days'	times	time's
tidig	early
tidiga	early
tidigare	earlier
tidigast	the earliest
tidigt	early
tidning	newspaper	journal
tidningar	magazines
tidningarna	papers
tidningen	the newspaper	paper
tidpunkt	date	time
tidpunkten	the time	the moment	time
tids	time
tidskrift	newspaper	magazine
tidskriften	the magazine
tidskrifter	magazines	periodicals
tidszon	timezone	time zone
tidszoner	time zones
tidvis	times
tiger	tiger	silent
tigern	the tiger
tigrar	tigers
till	to
tillbaka	back
tillbehör	condiments	accessory
tillbringade	spent
tillbringar	spends	spend
tilldelades	awarded
tilldelas	assigned	award
tilldelats	awarded
tillfälle	occasion	instance
tillfällen	occasion	oppertunities
tillfället	time
tillfällig	temporarily
tillfälliga	temporary
tillfälligt	temporarly	temporary
tillgänglig	available	provided
tillgängliga	available
tillgängligt	available
tillgång	access
tillgångar	assets
tillgången	access
tillhandahåller	provides
tillhör	belongs	belonging to
tillhöra	belong to	belonging to
tillhörande	belonging to	belonging (to)
tillhörde	was a part of	belonged to
tillhörighet	belonging	belonging; affiliation
tillhört	belonged	belonged to
tillika	also
tillkom	resided	hold back
tillkommer	reside
tillkommit	accured	been
tillkomst	origin	established	advent
tillkännagav	announced
tillräcklig	sufficient	enough
tillräckliga	insufficient	sufficient
tillräckligt	sufficient
tills	until the	until
tillsammans	together
tillstånd	to the dental	condition
tillståndet	condition	the state
tillsätts	appointed	appoints
tilltagande	increasing
tillträdde	assumed
tillträde	access
tillvaron	existence	the subsistence
tillverka	producing
tillverkade	manufactured	made
tillverkar	makes
tillverkare	producer	manufacturer
tillverkas	is made	manufacture
tillverkning	production
tillverkningen	production	the production
tillväxt	growth
tillväxten	growth
tilly	tilly
tillägg	addition
tillämpa	administer	implement	applying
tillämpar	administer	practice	administers
tillämpas	applied
tillämpningar	situations	implementations
tillät	distillate	allowed
tilläts	was allowed	allowed
tillåta	allow
tillåtelse	allowed	permission
tillåter	allows	allow
tillåtet	allowed
tillåtna	allowed
tillåts	is allowed	allowed
tim	h	tim
time	time
timmar	hours
timme	hour
tina	thaw	tina
ting	matters	thing
tingslag	leet
tintin	tintin
tio	ten
tionde	tenth
tiotusentals	tens of thousands
titanic	titanic
titanics	titanic's
titel	title
titeln	the title	title
titlar	titles
titta	watch
tittar	looking; viewing; viewer	viewing
tittarna	the viewers	viewers
tjeckien	czech republic	the czech republic
tjeckiska	czech
tjeckoslovakien	czechoslovakia
tjugo	twenty
tjäna	profit	make	earn
tjänade	earned
tjänar	earns	serves
tjänare	servant
tjänst	service
tjänstemän	officals	officials
tjänsten	service
tjänster	services
tobak	tobacco
tobias	tobias
tog	was	took
togs	taken	were taken
tokyo	tokyo
tolerans	tolerance
tolfte	twelth
tolka	interpreting	interpret
tolkade	interpreted
tolkar	interprets	views
tolkas	is interpreted	interpret
tolkats	interpret	interpreted
tolkien	tolkien
tolkiens	tolkien's
tolkning	interpretations	interpretation
tolkningar	interpretations	interpretation
tolkningen	interpretetation
tolv	twelve
tom	tom
tomas	tomas
tomma	empty
tomt	empty	blank
ton	tone
tongivande	influential
tony	tony
top	top
topp	top
toppade	topped
toppar	tops	(that) peaks
toppen	peak	the top
tor	thu	thor
torah	torah
torbjörn	torbjorn
torde	could
torg	square
torget	square	the square
torka	dry
torn	tower
tornen	towers	the tower
tornet	the tower
toronto	toronto
torra	dry
torres	torres
torrt	dry
torsten	torsten
tortyr	torture
tosh	tosh
total	total
totala	total
totalt	complete	wholly
tottenham	tottenham
tour	tour
toy	toy
tradition	tradition
traditionell	traditional
traditionella	traditional
traditionellt	traditional
traditionen	the tradition
traditioner	traditions	the traditions
traditionerna	traditions	the traditions
trafik	traffic
trafiken	traffic	the traffic
trafikerade	frequent
trafikerar	traffic	frequent
trafikeras	trafficked
trakten	the region	region	area
transeuropeiska	transeuropean
transkription	transcript
transport	transportation	transport
transporter	transports
transportera	transport
transporterar	transports
transporteras	is transported	transported
tre	three
tredje	third
tredjedel	a third
tredjedelar	thirds
tree	tree
treenigheten	tinity	the trinity
treenighetsläran	doctrine of the holy trinity	trinity	school of trinity
trend	trend
trenden	trend	the trend
trettio	thirty
trettioåriga	13 year olds	thirty year's (war)	thirty years
tretton	thirteen
trey	trey
triangel	triangle
triangeln	triangle	the triangle
triangelns	triangle	the triangle's
trianglar	traingles
trigonometriska	trigonometric
trinidad	trinidad
tro	believing	think
trodde	thought
troende	faithful
troligen	probably	likely
troligt	likely
troligtvis	probably
tron	faith
tronen	the throne
tronföljare	heir	successor
tropisk	tropical
tropiska	tropical	tropic
tropiskt	tropical
tror	believe	think
tros	belived
trosbekännelsen	creed
trossamfund	religious community	faith community
trots	although
trotskij	trotskij
truman	truman
trummis	drummer
trummisen	the drummer	drummer
trummor	drums
trupp	troops	troop
trupper	troops
trupperna	troops	the troops
tryck	print	pressure	press
trycket	pressure
tryckta	printed
trycktes	was published	printed
trä	wood
träd	into	tree
träda	emerge	fallow
trädde	come into effect	entered
träffa	meet	see
träffade	met
träffades	was met	reached; met
träffar	meets
träffas	meet	reached
träffat	met
tränade	trained
tränare	coach
tränaren	the coach
tränga	push (aside)	cut in
tränger	forces forward	cut in
träning	training	practice
trådlös	wireless
trött	tired
tsar	tsar	czar
tsaren	the czar	the tsar
tsunami	tsunami
tsunamier	tsunamis
tum	inch	inches
tung	heavy
tunga	heavy	tongue
tungt	heavy
tunisien	tunisia
tunn	thin
tunna	thin
tunnel	tunnel
tunnelbana	subway
tunnelbanan	subway; tube; underground	the subway
tunnlar	tunnels
tupac	tupac
tur	turn	tour
turism	tourism
turismen	tourism	the tourism
turister	tourists
turistmål	tourist destination	tourist attraction
turkar	turks
turkarna	turks	the turks
turkiet	turklet	turkey
turkiets	turkey's	turkeys
turkisk	turkish
turkiska	turkish
turner	tournament
turnera	tour
turnerade	toured
turneringen	the tournament
turné	tour
turnéer	tours
turnén	tour	tournament
tusen	thousands
tusentals	thousands
tv	tv
tvfilm	tv-movie	tv film
tvinga	force
tvingade	forced
tvingades	forced
tvingas	forced
tvingats	forced
tvister	conflicts	disputes
tvkanaler	tv channels
tvprogram	tv program	tv-show
tvserie	tv serial
tvserien	tv series	the tv show	television program
tvserier	tv-shows	tv shows	tv-series
tvskådespelare	tv actor
tvungen	forced	forced (to)
tvungna	forced	forced to
tvärtom	on the contrary	contrary to
två	two
tvåa	second
twilight	twilight
ty	for
tycker	thinks
tyckte	thought
tycktes	seemed
tyder	indicates
tydlig	clear	obvious
tydliga	clear	obvious
tydligt	clear	obvious
tyngre	heavier
typ	kind of	type
typen	the type	type
typer	types	characters
typerna	the types	types
typisk	typical
typiska	typical
typiskt	typically	typical
tysk	german
tyska	german
tyskar	germans
tyskarna	the german	the germans
tyske	german
tyskland	germany
tysklands	germany's	germanys
tyskt	german
tyst	silent	quiet
tyvärr	unfortunately
täcka	thank
täcker	attacks	covers
täcks	covered	covers
täckt	covered	coated
tämligen	rather	fairly
tänder	teeth
tänderna	teeh
tänka	think
tänkande	thinking
tänkandet	thinking	the way of thinking
tänkare	thinker
tänker	thinking
tänkt	supposed; intended	intended
tänkte	thought	was going to
tät	compact	frequent
täta	close
tätbefolkade	densely populated	populated
tätort	urban	conurbation
tätorten	conurbation
tätorter	urban	cities	conurbation
tätt	tight	tightly
tävla	compete
tävlade	competed
tävling	competition	contest
tävlingar	competitions	contests
tävlingen	competition	contest
tåg	rail	trains
tågen	the trains
tåget	train	the train
tål	stand	is resistant to
u+	u +
udda	odd
uefa	uefa
uefacupen	the uefa champions league	uefacupen
uganda	uganda
ugandas	of uganda
uggla	owl
ugglas	owl	ugglas
uk	uk
ukraina	ukraine
ukrainas	ukranian	ukraine's
ukrainska	ukrainian
ulf	ulf
ullevi	ullevi
ulrich	ulrich
ultraviolett	ultraviolet
umgänge	company	intercourse
und	und
undan	away (from)	escape
undantag	exception	except
undantaget	except
under	during	under
underart	subspecies
underarten	subspecies	sub species
underarter	sub-species	subspecies
undergång	doom	destruction
underhåll	support	allowance	entertainment
underhållning	entertainment
underjordiska	underground
underliggande	underlying
underlätta	ease	facilitate
underlättar	make it easier
underordnade	subordinates	subordinate
undersöka	study	research
undersökning	survey
undersökningar	surveys; investigations	studies	studies'
undersökte	investigated	examined
undertecknades	signed
underverk	wonder
undervisade	taught
undervisning	education
undervisningen	the education
undre	lower
undvika	prevent	avoid
undviker	avoids
unesco	unesco
unescos	unesco
ung	young
unga	young
ungar	babies	kids; offsprings; young
ungarna	the kids	kids	the young
ungdom	youth
ungdomar	youths	adolescents	the youth
unge	young	kid
ungefär	approx.; approximately	approximately
ungern	hungaria
ungerns	hungary	hungrarys
ungerska	hungarian
uniform	uniform
unik	unique
unika	unique
unikt	unique
union	union
unionen	union	the union
unionens	the union	the union's
universitet	university
universiteten	universities	the universities
universitetet	the university	university
universum	universe
universums	the universe's	universe's
uno	uno
up	up
upp	up
uppbyggd	structered	built-up
uppbyggnad	construction	structure
uppbyggt	structured
uppdelad	divided	split
uppdelade	divided
uppdelat	divided	split
uppdelning	division	partitioning	playback
uppdelningen	division	partitioning; sectionalization; division; split (-ting)
uppdrag	job	missions	mission
uppdraget	task; assignment	assignment
uppe	top	up	(on) top, up, above
uppehåll	residence	pause	hiatus
uppemot	almost
uppenbarelse	revelation	apparition
uppenbarelser	revelations
uppfann	invented
uppfanns	was invented	invented
uppfatta	apprehend	perceive
uppfattade	perceived	perceive
uppfattar	percieves	interpret
uppfattas	perceived	are regarded
uppfattning	understanding
uppfattningar	opinions	perceptions
uppfattningen	comprehension
uppfinnare	inventor
uppfinningar	inventions
uppfostran	upbringing
uppfylla	satisfy	fulfill	meet (requirements)
uppfyller	fulfills
uppföljare	sequel
uppförande	behavior
uppfördes	was constructed	constructed
uppgav	said
uppger	states	state
uppges	reported
uppgick	total	was
uppgift	task	data
uppgiften	the task
uppgifter	information	tasks
uppgifterna	data	the information
uppgörelse	agreement	deal
upphov	origin	source	rise
upphovsman	creator	author
upphovsrätt	rise knob	copyright
upphovsrätten	copyright
upphörde	ceased	expired
upphört	ceased
uppkallad	named
uppkom	arose
uppkommer	arises	resulting	arises; generated
uppkommit	arisen
uppkomst	onset	origin
uppkomsten	onset	origin
upplaga	edition
upplagan	edition
upplagor	editions	issues
uppleva	experience
upplevde	felt	experienced
upplevelse	experience
upplevelser	experiences
upplever	experience
upplysning	the enlightenment	enlightenment
upplysningen	the enlightenment
upplysningstiden	enlightenment	age of enlightenment
upplösning	resolution; dissolution	resolution
upplösningen	disbandment
upplöstes	dissolved
uppmanade	urged	encouraged
uppmaning	call; injunction	exhortation
uppmuntrade	encouragement	encouraged
uppmärksamhet	attention	attantion
uppmärksammad	noted, come to attention	noticed
uppmärksammade	observed	noted	noticed
uppmärksammades	attention	drew attention
uppmärksammat	noticed
uppnå	achieving	achieve
uppnådde	met	achieved
uppnår	achieve	reaches
uppnås	is achieved
uppnått	met	achieved
upprepade	repeated
uppror	uprising	rebellion
upproret	the upprising	revolt
upprustning	renovation
upprätta	establish	up
upprättade	established	prepared
upprättades	was established	establish
upprättandet	establishment
upprättas	established	establish
upprätthålla	maintain	keep up
upprätthåller	maintains	maintaining
uppsala	uppsala
uppskatta	appreciate
uppskattad	estimated	appreciated
uppskattade	estimated	appreciated
uppskattades	estimated	appreciated	was appreciated
uppskattar	estimates
uppskattas	is appreciated	appreciated
uppskattning	appreciation
uppskattningar	estimates
uppskattningsvis	approximately
uppslagsordet	entry word	lexical entry; word
uppslagsverk	encyklopedia
uppstod	developed	was
uppstå	develop
uppståndelse	resurrection
uppstår	occur
uppstått	arised	arisen
uppsving	boost
uppsättning	equipment
upptagen	busy	occupied
upptar	occupies
uppträda	appear	occur
uppträdande	performance	appearance	conduct
uppträdde	appeared	perform	occurred
uppträder	occur	performs	appears
upptäcka	discover
upptäcker	discoveries
upptäcks	detected	discoverd	is discovered
upptäckt	discovered	discovery
upptäckte	discovered	found
upptäckten	the discovery
upptäckter	discoveries	discovery
upptäcktes	discovered	(was) discovered
uppvisade	showed
uppvisar	shows
uppvärmning	heating	warming
uppvärmningen	the warm-up	the warmup
uppväxt	growing up
uppåt	up	upwards
ur	from	out
uralbergen	the ural mountains
uran	uranium
urin	urine
urskilja	distinguish	discern
ursprung	origin	root
ursprunget	origin	the origin
ursprungliga	original
ursprungligen	originally
ursprungsbefolkning	native population
ursprungsbefolkningen	the native population	indigenous people	indigenous population
ursäkt	excuse
uruguay	uruguay
urval	selection
usa	the usa	united states of america	usa
usama	osama	usama
usas	usa:s	u.s.
ut	out; up	out
utan	without
utanför	outside
utbildad	formed	educated
utbildade	educated
utbildning	education
utbildningen	education
utbredd	widespread
utbredda	widespread
utbredning	distribution	distrubution
utbrett	wide	widespread
utbrott	outbreak	outbreaks
utbröt	erupted	broke out
utbud	availibility
utbyggda	expanded	expand
utbyggnad	addition	development	expansion
utbyggt	develpoed	built	extended
utbyte	trade
utdelades	distributed
utdöda	extinct
ute	absent	out
uteslutande	exclusivly	only	exclusively
utformade	designed
utformning	layout	shape	formation
utformningen	the layout	layout
utfärdade	issued
utför	perform
utföra	perform	out
utföras	performed
utförd	completed	performed
utförda	made	performed
utfördes	carried out	was carried out	preformed
utförs	out	is done
utfört	done
utgavs	was published	published
utgick	started
utgifter	expenditure	expenses
utgiven	published
utgivna	issued	published
utgivningen	the publication	the release
utgjorde	made up	comprised; consisted of
utgjordes	make up	comprised; consisted
utgångspunkt	starting point	point of departure
utgår	deleted
utgåva	edition	issue
utgåvan	the edition	issue
utgåvor	issues
utgör	make up	constitutes
utgöra	compose	make up
utgörs	consists of	make up
utifrån	from the outside	from
utkanten	the outskirts	outskirts
utkom	issued	(was) issued
utkämpades	fought
utlandet	foreign land	abroad
utlopp	outflow	outlet
utländsk	foreign	foregin
utländska	foreign
utlänningar	foreigners
utlösa	trigger
utlösning	release	ejaculation	trigger
utlöste	triggered
utmed	along
utmärkande	distinguishing
utmärkelsen	award	the award
utmärkelser	commendations
utmärker	characterizes	characterized
utmärks	are characterized	characterized
utmärkt	excellently	excellent; superb; marked by; characterized by
utnyttja	use
utnyttjade	used
utnyttjar	using	uses
utnyttjas	utilized	used
utnämndes	was declared	appointed
utom	except
utomeuropeiska	non-european
utomlands	abroad
utomliggande	external; ex-territorial
utomstående	outside people; outsiders	outsider
utredning	study	investigation
utredningen	investigation	the investigation
utrikes	foreign
utrikesminister	minister of foreign affairs
utrikespolitik	foreign affairs	forgein policy
utrikespolitiken	the foreign policy
utrikespolitiska	foreign policy	foreign political
utropade	exclaimed	cried out
utropades	proclaimed	was proclaimed
utrotning	extinction	extermination
utrustning	equipment	gear
utrymme	space
utsatt	exposed
utsatta	exposed
utsattes	subjected	exposed
utse	appoint	name
utsedd	appointed
utseende	appearance
utser	chooses	appoints
utses	is appointed	designated	appointed
utskott	committee	organ
utsläpp	emissions
utspelar	takes place	set
utsträckning	extent
utställning	exhibition
utsätts	exposed
utsåg	declared
utsågs	was	appointed	was appointed
utsöndras	secrete	exudes
uttal	pronunciation
uttalade	commented; made a comment; spoke about	spoke
uttalande	statement
uttalanden	statements
uttalas	pronounced	be pronounced
uttalat	outspoken
uttalet	the pronounciation
uttryck	expression
uttrycka	express
uttrycker	express	expressing	express (-es)
uttrycket	the expression
uttryckligen	explicitly
uttryckt	expressed
uttryckte	expressed
utvalda	selected	selected; chosen
utveckla	develop	developing
utvecklad	developed
utvecklade	oral
utvecklades	(was) developed
utvecklandet	development
utvecklar	develops
utvecklas	development
utvecklat	developed	evolved
utvecklats	developed
utveckling	development
utvecklingen	development	the development
utvidgade	expanded
utvidgning	enlargement; expansion
utvinna	extract
utvinns	extracted
utvisning	penalty
utåt	outwardly	out
utökade	expanded	increased
utökat	extended
utöva	exercise
utövade	exercised
utövar	carrying	exercise
utövas	is practised	exercised
vacker	beautiful
vackra	beautiful	fine
vad	what
vaginalt	vaginal
vagn	wagon	carrige
vagnar	carts	wagons	carriges
val	election	choice
valborg	valborg
vald	elected	selected
valda	chosen
valde	crowned	chose
valdes	representatives'	selected	chosen; elected
valen	the elections	elections
valet	the election
valla	valla	herd
valley	valley
vallhund	herder	herding dog
valrörelsen	election campaign
valt	chosen
valuta	currency	exchange
valutan	currency
vampyr	vampire
vampyren	the vampire
vampyrer	vampires
van	van
vana	familiar	used
vandrar	wanders	migrates
vanföreställningar	delusions
vanlig	ordinary	common
vanliga	ordinary	regular	usual
vanligare	more common
vanligast	most usual	most common
vanligaste	frequent	most common
vanligen	usually
vanligt	usual
vanligtvis	usually
vann	won
vanns	(was) won
vapen	weapons	weapon
vapnen	the weapons
vapnet	the weapon	the weapon; escutheon; coat of arms; arms; badge
var	was
vara	be
varade	lasted
varandra	each other
varandras	each others	each other's
varar	lasts
varav	of which	which
vardagen	the weekday
vardagliga	ordinary	everyday
vardagligt	everyday
vardera	either	each
vare	either
varefter	whereafter
varelse	creature
varelser	creatures
varför	why
varg	wolf
vargar	wolves
vargen	the wolf
variant	variant	type	variety
varianten	version	variant
varianter	variants	diversities
varianterna	the diversities
variation	diversity
variationer	variations
variera	vary
varierade	varied
varierande	variable	varied	varying
varierar	varies	vary
varierat	varied
varifrån	from where; wherefrom
varit	has been	been
varje	each
varken	neither	either
varm	warm
varma	hot	warm
varmare	warmer
varmblod	warmblood
varmed	whereby
varmt	hot	warm
varna	varna
varnade	warned
varning	warning
varor	products
varpå	thereafter	whereupon	after which
vars	whose	who's
varsin	(one) each	opposite
vart	each
varuhus	warehouse	department store
varv	dockyard	shipbuilding
varvid	in which
vasa	vasa
vasaloppet	vasaloppet
vasas	vasas	vasa's
vatikanstaten	vatican city	the vatican	vatican
vatten	water
vattendrag	streams	watercourse
vattenkraft	water power	hydroelectric power
vattenånga	steam	water vapour
vattnet	water	the water
vattnets	the water's	the waters
vd	ceo
vecka	week
veckan	weeks	the week
veckor	weeks
veckorna	weeks
vegas	vegas
velat	wanted
vem	who
venedig	venice	venedig
venezuela	venezuela
venus	venus
verde	verde
verk	work	works
verka	seem	operate	appear
verkade	were active, worked, was active
verkan	effect
verkar	seems	operates
verkat	worked	acted
verken	plants	wroks
verket	plant; indeed	plant
verklig	real
verkliga	real
verkligen	real	the reality
verklighet	true	reality
verkligheten	reality
verksam	active	effective
verksamhet	work	activity
verksamheten	the work	activity
verksamheter	operations	businesses	activity
verksamma	active
verkställande	executive
verktyg	tool	tools
vers	verse
versaillesfreden	treaty of versailles
version	version
versionen	edition	the version
versioner	versions
vet	know
veta	know
vete	wheat
vetenskap	science
vetenskapen	the science	science
vetenskaplig	learn scientific	scientific
vetenskapliga	scientific
vetenskapligt	scientifically	scientific
vetenskapsmän	scientist	scientists
veto	veto	vetoe
vhs	vhs
vi	we
via	via	through
vice	vice
vicepresident	vice president
victor	victor
victoria	victoria
victoriasjön	victoria lake	lake victoria
vid	at	by	in
vida	broad	wide
vidare	moreover	further
video	video
videon	the video
vidsträckta	broad	wide; broad
vidta	take
vietnam	vietnam
vietnamesiska	vietnamese
vietnamkriget	the vietnam war	vietnam war
vietnams	vietnam's
viggo	viggo
vii	vii
vika	fold
viken	gulf
viking	viking
vikingar	vikings
vikingarna	the vikings
vikingatiden	the viking age
vikt	weight
vikten	importance
viktig	major	important
viktiga	important
viktigare	more important
viktigaste	most important
viktigt	important
viktor	viktor
vila	rest
vilar	rests
vilda	wild
vilhelm	vilhelm
vilja	will
viljan	will	te will
vilka	who; which; that	who
vilkas	whose
vilken	which
vilket	which
vill	will	want
villa	house	villa
ville	wanted (to)	wanted
villkor	conditions	condition
villkoren	the terms	conditions
villor	houses	villas
vimmerby	vimmerby
vin	whine	wine
vincent	vincent
vinci	vinci
vind	wind
vindar	winds
vinden	the wind	wind
vindkraft	wind power
vindkraftverk	wind turbine	wind power station
vingar	wings
vinkel	angle
vinkeln	angle	the angle
vinklar	angles
vinna	win
vinnare	winner
vinnaren	winner	the winner
vinner	gaining	win	wins
vinst	profit	win
vinsten	the win
vinster	profit
vinter	winter
vintergatan	milky way	the milky way
vinterkriget	the winter war
vintern	the winter	winter
vinterspelen	winter games
vintertid	winter-time
vintrar	winters
vintrarna	the winters	winters
virginia	virginia
virus	virus
viruset	virus
vis	wise	way
visa	see
visade	showed	showed; displayed
visades	showed
visar	shows
visas	is showed	shown
visat	shown
visats	shown	demonstrated
visby	visby
visdom	wisdom
vision	vision
visor	songs
viss	certain
vissa	some
visserligen	certainly	although
visst	specific	certain
visste	did
vista	vista
vistas	live	present
vistelse	visit	stay
vit	white
vita	white
vitryssland	belarus
vitt	white	widely
vittne	witness
vittnen	witnesses
vladimir	vladimir
vm	world championship
voddler	voddler
vojvodina	voyvodina	vojvodina
vojvodskap	voivodeship
vol	v
voltaire	voltaire
volvo	volvo
volym	volume
von	von
vore	would	were
vrida	twist	turn
vulkaner	volcanos	volcanoes
vulkaniska	vulcanic	volcanic
vulkanutbrott	vulcano eruption	volcanic eruption
vunnit	won
vuxen	adult
vuxit	grown
vuxna	adult
väckt	awaken	woken
väckte	awakened	aroused
väder	weather
vädret	the weather
väg	vague	way
vägar	roads
vägarna	paths	roads (roadways)
vägen	the road	road
väger	weighs	weight
vägg	wall
vägnät	network
vägnätet	road network
vägrade	refused
vägrar	refuses	refuse
väl	selecting	good
väldet	empire	violence	the rule
väldiga	immense	vast
väldigt	very
välfärd	wealth	welfare
välgörenhet	charity
välja	select
väljas	elected	choose
väljer	elects
väljs	elect
välkänd	well-known	well known
välkända	well known
välmående	well-being; affluent	prosperous
välstånd	prosperity
vän	van	friend
vända	turn	habituated
vände	turned
vänder	turn
vännen	the friend	friend
vänner	friendas	friends
vänskap	friendship
vänster	left
vänstern	western	left party
vänsterpartiet	leftist party	left-wing party	left wing party
vänstra	left-hand	left
vänt	turned
vänta	(have to) wait; expect	wait
väntade	expected; were waiting	waited
väntan	awaiting	waiting	wait
väntar	waiting	expect
väntas	expected
väntat	expected
väpnad	armed
väpnade	armed
värd	worth
värde	value
värdefulla	valueable	valuable	value
värden	values
värderingar	evaluations	values
värdet	the value
värld	world
världen	world	the world
världens	the world's	the world	the worlds
världsarv	world heritage
världsarvslista	world heritage list
världsbanken	world bank
världsdel	continent
världshälsoorganisationen	world health organization
världskrigen	the world wars
världskriget	world war
världskrigets	the world war's	world war
världsliga	worldly
världsrekord	world record
världsturné	world tour
värme	thermal
värmestrålningen	heat radiation
värmland	wermlandia
värmlands	varmlands	värmlands	hot countries
värnplikt	military service
värnpliktiga	conscripted
värre	worse
värsta	worst
värt	worth
värvade	recruited
väsen	entity
väsentligt	substantially	relevant
väska	bag	fluid	pan	suitcase
väst	west	the west
västbanken	the west bank	westbank
västberlin	west berlin
väster	west
västerbottens	västerbottens	västerbotten's
västergötland	västergötland
västerländsk	western
västerländska	western
västerut	westward; west	westwards
västerås	västerås
västeuropa	western europe
västindien	west india
västkusten	the west coast
västlig	western
västliga	western
västmakterna	western powers
västra	west	vastra	western
västsahara	western sahara
västtyskland	west germany
västvärlden	western world
väte	hydrogen
vätet	the hydrogen
vätska	fluid
växa	grow	wax
växande	growing
växer	grows
växjö	växjö
växt	plant
växte	grew
växter	plants
växterna	plants
växthuseffekten	the greenhouse effect
växthusgaser	vaxthusgaser	greenhouse gas
våg	vague	road	wave
vågade	dared
vågen	the wave
våglängder	wavelengths	wave lengths
vågor	waves
våld	violence
våldet	the violence	violence
våldsam	violent
våldsamma	violent
våningar	floors	storeys
vår	spring
våra	our
vård	vard	nursing	healthcare
våren	spring	the spring
vårt	our	each
w	w
wagner	wagner
wahlgren	wahlgren
wailers	wailers
wales	wales
wall	wall
wallace	wallace
wallander	wallander
wallenberg	wallenberg
wallenstein	wallenstein
walt	walt
walter	walter
want	want
war	war
warhol	warhol
warner	warner
warszawa	warzaw	warsaw
washington	washington
waterloo	waterlo	waterloo
watson	watson
way	väg
wayne	wayne
we	we
webbkällor	websources	web sources
webbplats	website
webbplatsen	webpage	the website	site
webbplatser	webbsites	websites
weber	weber
welsh	welsh
wembley	wembley
werner	werner
west	west
what	what
who	who
wien	vienna
wikipedia	wikipedia
wikipedias	wikipedias
wild	wild
wilde	wilde
wilhelm	wilhelm
will	will
william	william
williams	williams
willy	willy
wilson	wilson
wind	wind
winnerbäck	winnerbäck	winnerback
winston	winston
without	without
wittenberg	wittenberg
wolfgang	wolfgang
works	works
world	world
wright	wright
x	x
xi	xi
xii	xii
xiis	xii
xis	the eleventh's
yngre	younger
yngsta	youngest
yngste	youngest
york	york
yorks	yorks
you	you
youtube	youtube
yta	surface
ytan	the area	surface	area
ytterligare	further	additional
ytterst	very; extremely	highly
yttersta	furthest	supreme	highly
yttre	outer
z	z
zach	zach
zagreb	capital of croatia	zagreb
zanzibar	zanzibar
zarathustra	zarathustra
zeeland	zeeland
zeppelin	zeppelin
zeus	zeus
zink	zinc
zirkon	zirkon	zirconium	zircon
zlatan	zlatan
zon	zone
zonen	the zone	zone
zoner	zones
zuckerberg	zuckerberg
 cm	centimeters	cm
 kilometer	kilometer
 km	kilometers
 kmh	km/h
 km²	kilometres
 meter	metre	meter
 miljoner	millon	one million	millions
 mm	millimeter
 procent	percent	per
  km²	square kilometre	km²	km2
 °c	celsius
£m	million pounds
×	x
à	river
äga	own	aga
ägande	owning
ägare	owner
ägda	owned
ägde	tookplace; occured	owned
ägdes	owned
äger	owns
ägg	egg
ägna	spend	devote
ägnade	dedicated
ägnar	spend time	dedicated	spends time
ägs	is owned	(is) owned
ägt	taken
äkta	married	genuine
äktenskap	the marriage	marriage
äktenskapet	marriage
äldre	older
äldsta	oldest
äldste	elders	eldest
älg	moose
älgar	moose
älgen	elk; moose
älska	love
älskade	loved	loved; beloved
älskar	loves
ämbetsmän	officers	bailies	officer
ämne	substance
ämnen	agents
ämnena	subjects	the elements	substances
ämnet	substance	subject
än	yet	than
ända	as far as
ändamål	purpose
ände	end
änden	end	spirit
ändra	change
ändrade	changed
ändrades	changed	was
ändrar	changing	changes
ändras	be changed
ändrat	changed
ändringar	edit	changes
ändå	still	spirit
änglar	angels
ängssyra	sorrels	sorrel	sorell
ännu	still	yet
är	is
ära	oar	glory
ärftliga	genetic
ärkebiskop	archbishop
ärkebiskopen	archbishop
äta	eat
äter	eats	eat
ätten	the dynasty
ättlingar	descendants
även	also
äventyr	adventure	adventures
å	on	river
åka	go
åke	åke
åker	go	field; going
åkte	went	relegated
åland	Åland
ålands	Åland island's	the Åland island's
ålder	age
åländska	Åland swedish
ån	on	the river
ångest	anxiety	anguish
år	the year	year
åren	the years	years
årens	the year's	years
året	all year	the year
årets	the year's
århundraden	centuries
århundradena	centuries
århundradet	century
årig	year old
åriga	-year	year
åring	year old	years
årlig	yearly
årliga	annual
årligen	annually	yearly
års	years (age)	years
årsdag	anniversary
årstiderna	the seasons
årsåldern	age group	years old
årtionde	decade
årtionden	decades
ås	ridge
åsikt	opinion
åsikten	the opinion	view
åsikter	opinions
åskådare	spectators	audience; viewer
åstadkomma	provide	create
åt	to	for
åtal	prosecution
åtalades	was prosecuted	charged
åter	again
återfanns	was rediscovered	can be found
återfinns	is rediscovered
återförening	reunion
återgick	returned	returning
återigen	once again	yet again
återkom	return	feedback	returned
återkommande	recurring
återkommer	returning
återkomst	return
återställa	resett
återstående	remaining
återstår	remains	remain
återta	regain	retake	reclaim
återvända	return
återvände	returned	returning
återvänder	returns	atervander
återvänt	returned
åtgärder	measures
åtminstone	at least
åtskilda	segregated	separate
åtskilliga	several
åtta	eight
åttonde	the eighth
ö	o
öar	islands
öarna	the islands	islands
öde	fate
ödleblad	lizardtail	ödleblad	lizard blade	houttuynia cordata	odleblad	lizardleaf	lizard tail	chameleon plant
öga	eye
ögat	eye
ögon	eye (-s)	eyes
ögonen	eyes
öka	oka	increase
ökad	increase	increased
ökade	increased
ökande	increasing	rising
ökar	increases
ökat	increased
öken	desert
ökenråttor	gerbil	desert rats	gherbils	okenrattor	gerbils; desert rats	gerbils
öknen	the desert	desert
ökning	increase
ökningen	increase	the increase
öl	beer
öland	oland	öland
ölet	the beer	beer
ön	island	the island
öns	the islands	island's
önskade	desired	wished
önskan	desired
önskar	wish	desired
önskemål	desire	requests	demands
öppen	open
öppet	open
öppna	open
öppnade	opened	opening
öppnades	were opened	was opened	opened
öppnat	opened
örebro	Örebro
öresund	the sound
öron	ears
öronen	the ears
öst	east
östafrika	east africa
östasien	east asia
östberg	Östberg
östberlin	east berlin
östblocket	east block	the eastern bloc	cheese block
öster	east
östergötland	Östergötland
österrike	austria
österrikes	austria's	austrias
österrikeungern	oster kingdom hungary	austria-hungary
österrikiska	austrian
östersjön	baltic	balticsea
österut	eastwards	east
östeuropa	eastern europe	east europe
östfronten	eastern front	the east front
östman	Östman
östra	eastern
östtimor	east timor
östtyska	east german
östtyskland	east germany
östtysklands	east germany's	osttysklands
över	over
överallt	everywhere	overall; everywhere
överbefälhavare	commander-in-chief
överens	in agreement	agree
överenskommelse	deal
överensstämmer	conform	agree
överföra	transmit	transfer
överföras	transfer	transferred
överföring	transfer
överförs	is transferred	transfered
övergav	abandoned
övergick	transended	went over	switched
övergrepp	assult (-s)	abuse	assault
övergripande	over arching	general
övergå	transition	transend
övergång	transition
övergången	the transition	transformation
övergår	surpasses	released	exceed
överhuvudtaget	on the whole
överhöghet	suzeranity	supremacy	sovereignty
överleva	survive
överlevande	survivor; survivors; surviving
överlevde	survived
överlever	survives
överlevnad	survival
överlevt	survived
överlägset	superior
övernaturliga	supernatural	over natural
överraskande	surprisingly
övers	transl	translation
översatt	translated
översikt	overview	over term
överst	at the top; uppermost
översvämningar	floodings
översättas	translated	be translated	translated (to)
översättning	translation
översättningar	translations
översättningen	the translation
översätts	translate	is translated
övertala	convince	persuade
övertalade	over spoke	persuaded
övertog	took over	overtook
övertogs	overtaken
övertyga	convince
övervikt	obesity	overweight
övervägande	the predominant	predominant
övre	upper
övrig	other
övriga	other	others
övrigt	other
